��b   ˀ� ��                                                                            �                                                                                                                                                                                                                            @                  ��                                                                            �                                                                                                                                                                                                                            @                  ��                                                                            �                                                                                                                                                                                                                            @                  ��                                                                            �                                                                                                                                                                                                                            @                  ��                                                                           �                    ����������������������������������������                                                                                                                                                               @                  ��                  ���������������������������������������                  �                    �                                                                                                                                                                                                      @                  ��                  ���������������������������������������                  �                    �                                                                                                                                                                                                      @                  ��                  ���������������������������������������                  �                    �                                                                                                                                                                                                      @                  ��                  ���������������������������������������                  �                    �                                                                                                                                                                                                      @                  ��                  ���������������������������������������                  �                    �                                                                                                                                                                                                      @                  ��                  ���������������������������������������                  �                    �                                                                                                                                                                                                      @                  ��                  ���������������������������������������                  �                    �                                                                                                                                                                                                      @                  ��                  ���������������������������������������                  �                    �                                                                                                                                                                                                      @                  ��                  ���������������������������������������                  �                    �                                                                                                                                                                                                      @                  ��                  ���������������������������������������                  �                    �                                                                                                                                                                                                      @                  ��                  ���������������������������������������                  �                    �                                                                                                                                                                                                      @                  ��                  ���������������������������������������                  �                    �                                                                                                                                                                                                      @                  ��                  ���������������������������������������                  �                    �                                                                                                                                                                                                      @                  ��                  ���������������������������������������                  �                    �                                                                                                                                                                                                      @                  ��                  ���������������������������������������                  �                    �                                                                                                                                                                                                      @                  ��                  ���������������������������������������                  �                    �                                                                                                                                                                                                      @                  ��                  ���������������������������������������                  �                    �                                                                                                                                                                                                      @                  ��                  ���������������������������������������                  �                    �                                                                                                                                                                                                      @                  ��                  ���������������������������������������                  �                    �                                                                                                                                                                                                      @                  ��                  ���������������������������������������                  �                    �                                                                                                                                                                                                      @                  ��                  ���������������������������������������                  �                    �                                                                                                                                                                                                      @                  ��                  ���������������������������������������                  �                    �                                                                                                                                                                                                      @                  ��                 ��������������������������������������� @                �                    �                                                                                                                                                                                                      @                  ��                 ��������������������������������������� @                �                    �                                                                                                                                                                                                      @                  ��                 ��������������������������������������� @                �                    �                                                                                                                                                                                                      @                  ��                 ��������������������������������������� @                �                    �                                                                                                                                                                                                      @                  ��                 ��������������������������������������� @                �                    �                                                                                                                                                                                                      @                  ��                 ��������������������������������������� @                �                    �                                                                                                                                                                                                      @                  ��                 ��������������������������������������� @                �                    �                                                                                                                                                                                                      @                  ��                 ��������������������������������������� @                �                    �                                                                                                                                                                                                      @                  ��                 ��������������������������������������� @                �                    �                                                                                                                                                                                                      @                  ��                 ��������������������������������������� @                �                    �                                                                                                                                                                                                      @                  ��                 ��������������������������������������� @                �                    �                                                                                                                                                                                                      @                  ��                 ��������������������������������������� @                �                    �                                                                                                                                                                                                      @                  ��                 ��������������������������������������� @                �                    �                                                                                                                                                                                                      @                  ��                 ��������������������������������������� @                �                    �                                                                                                                                                                                                      @                  ��                 ��������������������������������������� @                �                    �                                                                                                                                                                                                      @                  ��                 ��������������������������������������� @                �                    �                                                                                                                                                                                                      @                  ��                 ��������������������������������������� @                �                    �                                                                                                                                                                                                      @                  ��                 ��������������������������������������� @                �                    �                                                                                                                                                                                                      @                  ��                 ��������������������������������������� @                �                    �                                                                                                                                                                                                      @                  ��                 ��������������������������������������� @                �                    �                                                                                                                                                                                                      @                  ��                 ��������������������������������������� @                �                    �                                                                                                                                                                                                      @                  ��                 ��������������������������������������� @                �                    �                                                                                                                                                                                                      @                  ��                 ��������������������������������������� @                �                    �                                                                                                                                                                                                      @                  ��                 ��������������������������������������� @                �                    �                                                                                                                                                                                                      @                  ��                 ��������������������������������?������ @                �                    �                                �                                                                               �                                                                             �       @                  ��                 �������������������������������������� @                �                    �                               �                                                                              �                                                                            �       @                  ��                 �������������������������������������� @                �                    �                               �                                                                              �                                                                            �       @                  ��                 �������������������������������������� @                �                    �                               �                                                                              �                                                                            �       @                  ��                 �������������������������������������� @                �                    �                               �                                                                              �                                                                            �       @                  ��                 �������������������������������������� @                �                    �                              �                                                                             �                                                                           �       @                  ��                 ���������?���������������������������� @                �                    �         �                    ?�                                                        �                    ?�                                                      �                    ?�       @                  ��                 ������������������������������������� @                �                    �        �                    �                                                       �                    �                                                     �                    �       @                  ��                 ������������������������������������� @                �                    �        � ~                   �                                                       � ~                   �                                                     � ~                   �       @                  ��                  ������������������������������������                  �                   �       ��                   �       @                                              ��                   �                                                    ��                   �       @                  ��                  �����������������������������������                  �                   �       ��                   �       @                                              ��                   �                                                    ��                   �       @                  ��                  �������� ���������������������������                  �                   �       ?���                   �       @                                              ?���                   �                                                    ?���                   �       @                  ��                  �������� ���������������������������                  �                   �       ���                   �       @                                              ���                   �                                                    ���                   �       @                  ��                  �������  ���������������������������                  �                   �      ����                   �       @                                             ����                   �                                                   ����                   �       @                  ��                  ������� p���������������������������                  �                   �      ����                   ?�       @                                             ����                   ?�                                                   ����                   ?�       @                  ��                  ���������������������������������������                  �                   �                                        @                                             ���                   ?�                                                   ���                   ?�       @                  ��                  ���������������������������������������                  �                   �                                        @                                             ���                   ?�                                                   ���                   ?�       @                  ��                  ���������������������������������������                  �                   �                                        @                                             ���       �  `        �                                                   ���       �  `        �       @                  ��                  ���������������������������������������                  �                   �                                        @                                             ?���       �  |        o�                                                   ?���       �  |        o�       @                  ��                  ���������������������������������������                  �                   �                                        @                                             ���      a� 0�   `    o�                                                   ���      a� 0�   `    o�       @                  ��                  ���������������������������������������                  �                   �                                        @                                             �� ���   �� |�  �   �                                                   �� ���   �� |�  �   �       @                  ��                  ���������������������������������������                  �                   �                                        @                                            �� p��  ��� ��  � �o�                                                  �� p��  ��� ��  � �o�       @                  ��                  ���������������������������������������                  �                   �                                        @                                            �  p�� ?��� ��  � ?�<�                                                  �  p�� ?��� ��  � ?�<�       @                  ��                  ���������������������������������������                  �                   �                                        @                                            �  `�� >�����  �� ��                                                  �  `�� >�����  �� ��       @                  ��                  ���������������������������������������                  �                   �                                        @                                            �  ��� ������� ����                                                   �  ��� ������� ����        @                  ��                  ���������?�� 8 � ��`����������                  �                   �                                        @                                            � ���������� ����                                                   � ���������� ����        @                  ��                  ���������� ��< � �������������                  �                   �                                        @                                            �   ��������� ?���                                                   �   ��������� ?���        @                  ��                  ����������~ �?�> � �������������                  �                   �                                        @                                            �   ���?���� �� ���                                                   �   ���?���� �� ���        @                  ��                  ����������� �?�< � ���?����������                  �                   �                                        @                                            7�   �������� ~���                                                   7�   �������� ~���        @                  ��                  ����������� ��|��` ��?��?��������                  �                   �                                        @                                            ?�   ?����?��� ���?�                                                   ?�   ?����?��� ���?�        @                  ��                  ����������� ?��|� �` ~�?����������                  �                   �                                        @                                            o�   ?���?�?��������                                                   o�   ?���?�?��������        @                  ��                  ������?����� ? ��|� ~@ >�����������                  �                   �                                        @                                            �   >��� ����������                                                    �   >��� ����������         @                  ��                  ����� ?����� ? ��y� |� >��?���������                  �                   �                                        @                                            ��   ~}��� ���?������                                                    ��   ~}��� ���?������         @                  ��                  ����� ���� >���� |� <������������                  �                   �                                        @                                            ��   ~���� y��<���{ �                                                    ��   ~���� y��<���{ �         @                  ��                  ���������� ~��� <�� ������������                  �                   �                                        @                                            �   ���� ?���|��� ?�                                                     �   ���� ?���|��� ?�          @                  ��                  ���������������������������������������                  �                   �     ?    ����� ~��|?�� ?�          @                                                                                                                          ?    ����� ~��|?�� ?�          @                  ��                  ���������������������������������������                  �                   �     ?    ����� ~�?�����  8        @                                                                                                                          ?    ����� ~�?�����  8        @                  ��                  ���������������������������������������                  �                   �     ?   ������ �������  0        @                                                                                                                          ?   ������ �������  0        @                  ��                  ���������������������������������������                  �                   �       ������ 8������  0        @                                                                                                                            ������ 8������  0        @                  ��                  ���������������������������������������                  �                   �       ?� �� x����� |�  0        @                                                                                                                            ?� �� x����� |�  0        @                  ��                  ���������������������������������������                  �                   �      �� �������� �?�           @                                                                                                                           �� �������� �?�           @                  ��                  ���������������������������������������                  �           ������� �     ? �� �������?�  �        G�������                                                                                                                   ? �� �������?�  �        @                  ��                 ��������������������������������������� @                �          �������� �     ? �� �����~�?��?� �        G�������                                                                                                                   ? �� �����~�?��?� �        @                  ��                 ��������������������������������������� @                �          �������� �     ?��� ������~��� ��       G��������                                                                                                                  ?��� ������~��� ��       @                  ��                 ��������������������������������������� @                �          �������� �     ���� �� ?������� ��       G��������                                                                                                                  ���� �� ?������� ��       @                  ��                 ������ ���� ��8�� !���� ������ @                �         ��������� �     ���� >�� ?������ � ��       G��������                                                                                                                  ���� >�� ?������ � ��       @                  ��                 ������ ��?��� ��0��O� ����� ������� @                �         ��������� �     �� � ~�� ?�`��� ?  �        G���������                                                                                                                 �� � ~�� ?�`��� ?  �        @                  ��                 ������ ��?��� ���c��1�� ����� ������ @                �         ?��������� �      �� � < �  � ?� ��   ��       G���������                                                                                                                  �� � < �  � ?� ��   ��       @                  ��                 ����������������������������� ������ @                �        ���������� �              � ?�      ��       G���������                                                                                                                          � ?�      ��       @                  ��                 ����������������� ��?����������?������ @                �        ���������� �               �� �        �       G����������                                                                                                                          �� �        �       @                  ��                 ����������������� ��?����������������� @                �        ?���������� �                �� �                 G����������                                                                                                                           �� �                 @                  ��                 ����������������� ������������������� @                �        ����������� �                �  �         �       G����������                                                                                                                           �  �         �       @                  ��                 ����������������� �������������������� @                �       ����������� �                 �  �                  G�����������                                                                                                                           �  �                  @                  ��                 ����������������� �������������������� @                �       ����������� �                 �  �                  G�����������                                                                                                                           �  �                  @                  ��                 ����������������� �������������������� @                �       ������������ �                 �  �                  G�����������                                                                                                                           �  �                  @                  ��                 ��������������������������������������� @                �      ������������ �                                        G�����������                                                                                                                           �  �                  @                  ��                 ��������������������������������������� @                �      ������������ �                                        G������������                                                                                                                          �                     @                  ��                 ��������������������������������������� @                �      ������������ �                                        G������������                                                                                                                          >                     @                  ��                 ��������������������������������������� @                �     ������������� �                                        G������������                                                                                                                          >                     @                  ��                 ��������������������������������������� @                �     ������������� �                                        G�������������                                                                                                                                              @                  ��                 ��������������������������������������� @                �     ������������� �                                        G�������������                                                                                                                                              @                  ��                 ��������������������������������������� @                �    �������������� �                                        G�������������                                                                                                                         8                     @                  ��                 ��������������������������������������� @                �    �������������� �                                        G��������������                                                                                                                        0                     @                  ��                 ��������������������������������������� @                �    ?�������������� �                                        G��������������                                                                                                                        0                     @                  ��                 ��������������������������������������� @                �   ��������������� �                                        G��������������                                                                                                                        0                     @                  ��                 ��������������������������������������� @                �   ��������������� �                                        G���������������                                                                                                                                              @                  ��                 ��������������������������������������� @                �   ?��������������� �                                        G���������������                                                                                                                                              @                  ��                 ��������������������������������������� @                �   ���������������� �                                        G���������������                                                                                                                                              @                  ��                 ��������������������������������������� @                �  ���������������� �                                        G����������������                                                                                                                                             @                  ��                 ��������������������������������������� @                �  ���������������� �                                        G����������������                                                                                                                                             @                  ��                 ��������������������������������������� @                �                   �                                        @                                                                                                                                                             @                  ��                 ��������������������������������������� @                �                   �                                        @                                                                                                                                                             @                  ��                 ��������������������������������������� @                �                   �                                        @                                                                                                                                                             @                  ��                 ��������������������������������������� @                �                   �          � �   `� `               @                                                 � �   `� `                                                               � �   `� `               @                  ��                 ��������������������������������������� @                �                   �           � �        0             @                                                  � �        0                                                              � �        0             @                  ��                  ���������������������������������������                  �                    �           � �        0                                                               � �        0            @                                                 � �        0             @                  ��                  ���������������������������������������                  �                    �           ������ �g��g�8                                                              ������ �g��g�8            @                 p                               ������ �g��g�8             @                  ��                  ���������������������������������������                  ������������������ �           �`͛6��l��3lٰ             �����������������p                              �`͛6��l��3lٰ            @                 �                               �`͛6��l��3lٰ             @                  ������������������� ��������������������������������������� ������������������                   �           �`��6��l3o�0                               �*�                             �`��6��l3o�0            @                T                               �`��6��l3o�0             @                  ������������������� �����������9�2|�3�|����̓�������������� ������������������                   �                                                          �$�                             �`̓6��l3l0            @                $                                                            @                  ������������������� �����������9�2d�3�d�$��̓&O������������ ������������������                   �                                                          �(�                             �`͛6��l�3lٰ            @                D                                                            @                  ������������������� �����������<?	3?�f|��p������������ ������������������                   �                                                          p                              ��������g��g�l           @                 �                                                            @                  ������������������� �������������������������������������� ������������������                    �                                                           �����������������                 0�      `              G�����������������p                                                            @                  ��                  ��������������������������������������                  �                    �                                                                                             �        `              @                                                                              @                  ��                  ���������������������������������������                  �                    �                                                                                                                      @                                                                              @                  ��                  ���������������������������������������                  �                    �                                                                                                                      @                                                                              @                  ��                  ���������������������������������������                  �                    �                                                                                                                      @                                                                              @                  ��                  ���������������������������������������                  �                    �                                                                                                                      @                                                                              @                  ��                  ���������������������������������������                  �                    �                                                                                                                      @                                                                              @                  ��                  ���������������������������������������                  �                    �                                                                                                                      @                                                                              @                  ��                  ���������������������������������������                  �                    �                                                                                                                      @                                                                              @                  ��                  ���������������������������������������                  �                    �                                                                                                                      @                                                                              @                  ��                  ���������������������������������������                  �                    �                                                                                                                      @                                                                              @                  ��                  ���������������������������������������                  �                    �                                                                                                                      @                                                                              @                  ��                  ���������������������������������������                  �                    �                                                                                                                      @                                                                              @                  ��                  ���������������������������������������                  �                    �                                                                                                                      @                                                                              @                  ��                  ���������������������������������������                  �                    �                                                                                                                      @                                                                              @                  ��                  ���������������������������������������                  �                    �                                                                                                                      @                                                                              @                  ��                  ���������������������������������������                  �                    �                                                                                                                      @                                                                              @                  ��                  ���������������������������������������                  �                    �                                                                                                                      @                                                                              @                  ��                  ���������������������������������������                  �                    �                                                                                                                      @                                                                              @                  ��                  ���������������������������������������                  �                    �                                                                                                                      @                                                                              @                  ��                  ���������������������������������������                  �                    �                                                                                                                      @                                                                              @                  ��                  ���������������������������������������                  �                    �                                                                                                                      @                                                                              @                  ��                  ���������������������������������������                  �                    �                                                                                                                      @                                                                              @                  ��                  ���������������������������������������                  �                    �                                                                                                                      @                                                                              @                  ��                  ���������������������������������������                  �                    �                                                                                                                      @                                                                              @                  ��                  ���������������������������������������                  �                    �                                                                                                                      @                                                                              @                  ��                 ��������������������������������������� @                �                    �                                                                                                                      @                                                                              @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              