�)X        x   �   �   �   �       �   �   �   �   x                                                                                                           x               x   �   �   �   �   x                                     x               x               x                                         �   �   �   �   x                                                     x   �   �   �   �   x               x                                     x   �   �   �   �   x   �   �   �   �   x                                     x                                                                     x   �   �   �   �   x   �   �   �   �   x                                     x   �   �   �   �   x               x                                