��d  ��Q Q  g�����0   �    �                         �������   @ ?�                        ����d   ��� �      ?�                 n��?���    ?� D    ��                �������   c���                      ���  <���  H����	     `                 _�t  /�`  �t  0�  �   �             ���   ���  @�  �       0 @            ��   >1��  g   ��    ��    �            �\@ �<��  �@ �= P   #�  ��         �    ��� ��� �� ��   G  ��       �    /�a  �?� q  �  �  ���       �    [��  >@q�� $�  >`��    ?�       >     ��  y ���(	�  y��
 @  ~ 0     x     ��, � w��@. � p  �  �    �     o� ��  ;� �& ��  8� 8 ��� L     ��    _���� 7� �l\��� 6� 8���     ���   ��x��� �� X|���  @ 8���     8���   ��x?��� ��@�x?��� �  @0?���    0?���    ~ x?��� ?��0�?��� @  �p������   p?���    @p�������`������  �q������   p���� � ��p?�z����?�z��   s�w�� �   p?$r�   ��p����������`  w�p� �   pp� @ ��p� � ��������� �  �p� `   p� �   � p�� �� ��������� �  �� �� `   p�� ��   � x�L�� W� x��� X  ���� 0   x�@��  � |����� _� |��3��X  ���� 0   |�����  � �� ���k� ������l  �  �    �  _�  � ������+� ������,  �� ���   �� ��� � ��� ���/� �������,  �����   ?�� ��� � �������� ������  ?������   ?� ��� � ߟ������, ߟ�!���  ?�=���   �  |�� ���~���,￀ ���  ��?��   �  >�� ��>�>��,�? ~�  ��ߟ�ό   <  � ��z@�/~ Z�\�z�b��[   �^�_ǆ   x  ~  �������
�\���P��   z��~#�    � x  ����7��\�7�    �����!�      0  �����/��\�X/�    ����� �          ��s���^���    �_�w� �     �    ��(�
���^�"��    ����� v          ��X��K�^�"�K    ����� 6          ��(�
��_�"�    ����� 6          ��S��+�^���+ !  �_�w�      �    ���ǈ�+�_�	H�+  � �����           �������_���  @����           �����п��[���P��   z��             ���zs��?����������  }\_      x O   ����.��-�� .� }����    <     ���~���,���  �� �>���p   �>  >   �>߁����,~߂ �� �?}�~       |   ��������?���c��   ���     � �   �������+�������(   ���     ��   ��?���� /��������,   ��     ��   � <9���~ /� �������h   C���     ���   �  ~��� W� ?��� P   ���� �8     ��   �  �?� _� ���@X   � ��0     >�    � ����� �����t��@�    �  �p     p     � ����� ��������@�       �`            ��������_��������@         �          @ �������� �������`         �          @ `����ǂ���`����ǂ�  �      �          � p �������p �������  �     �         � �� ?������@� ?�����  `                 �� ����� L ����  0                 �� ����� 6 ���                   ��  o�� � ���l                   ���  _��� /� �       (           ���   ���@� _  ?�        p         0  �t>  ?�  w�>  ?`   � �   �         `  =����  ~�� ���  ~�   ��   �   ��    �  ����  ��  ���  �    p    �    @       ���� ���   w�� �     8         0       ��  ��x  �9�  � �       <            ��@  7��  p  4 @   �   �         0   ���  ���  �  |�    �  �     �   �   ��c��_��   c��`      �  �      `       ���?���    \?��     ?��              }������    ��       ���       ��     �������      ���        �         ?�      �������   @ �                          �������                                                                   Q Q  g�����0   �    �                         �������   @                           �����d   �     �                         n�������         D                        �������    �                         ��������  H �� 	      �                _�����`  � � �   ��              ��������  @ q���       8  @            ���  8���  ����    � p    �            ��0 �?��  > �  P   �  �         @    ��� ���  � �      ��       �    /��  <'��  � ><$     ��             [��  <�3�� $ a� |��      ?         <     ��R  z 	���( �  � 9 
 @ ,  |        x     ��� � ���@� � �  \ �      �     o�L �� ?� �L ��  � � ����     ��     _�����?� ����� � 8��� �    ���    ��X��� ��� ���� � @0��� `    ���    ��X?��� O��@X?��� H   0?��� 0   ?���    �0?��� ����?��� D   p�����8    0?���    �0����!���$�����"   q�����    0����   ���?�z��� l�?�z��   s�w��    p?$r�  ������	�� X�����	    w�p�    pp�   �p� �� �p������  `��p�    p� �   ��p�� ���� �p������  @��� ��    p�� ��  �@x�L����@x����  �������   x�@�� � �@��������`���3���  ������   |����� � �@�� ����`������B�  ��  ���   �  _� � ��?������_���������`  �� ����   ?�� ���@ ����� ������������`  ������   ?�� ���@ ���������/� �������0  ?�������   ?� ���  � ߟ��������ߟ�!����  ?�=���`   �  |��  ���~���￀ ���  ��?��`   �  >��  ��>�>п���? ~�  ��ߟ��`   <  �  ��z@�/~ ����z�b���  �^�_�`   x  ~   �������W����P��X  z��~#�    � x  ����7�W��7�X   �����!�      0  �����/�_��X/�X   ����� �          ��s��_����X   �_�w� �     �    ��(�
�߀�"��   ����� 0          ��X��߀��"��   ����� 0          ��(�
�[���"��   ����� 0          ��S��[����\ � �_�w� 0     �    ���ǈ�[�C�	H�\ � ����� 0          �����_����X @���� 0          �����п�_����P��X  z��  0           �a�zs��?������������ }\_  p    x O    �y��.����� .�� }���� p  <      �?��~�������  ��� �>���p `  �>  >    �߁��瀿��߂ �瀰 �?}�~ `      |    ��������/�����c��0   ��� �    � �    ��������_��������@   ��� �    ��  @ ���?�������������`   �� �    ��  @ �@<9���~��`��������  � C����    ���  � �@ ~�����`?����  � ���� ��     ��  � �` �?���p���D�  � � ���     >�   � �����������t��E   @  �  ��     p    �������	�� ������I�  @     �            �X������� ������ʀ                     ��������� L������   0                  �����Ǧ���&����ǧ                     � �������3 ������                    ��?���W��@�?����        8           ��������� 
�����       p            ��@���_�� @���P   �    �         @  ��� ��� � ����   �   �    �     �  ��X  ��X /� =@   �   �    @       ��$   2���@ � _  r�   x                 �� >  e��   S>  �     <��              =���� ���  �� �     ?   |     8      ��� '��  
� $    �   �             ���� 8���   �� 8�     �  �     �   �   �q��_�x  � q��` �    �  ?�      p      �������   ,�  @    ��             ��������   ��      ���       ��    ���������    ���        �         �      ���������     �                           }�������                                   �������                                    �������   @                             �������                                                                   Q Q  g�����0   �8  �                         �?���}�   @�  �                      ~�����d   �    @�                        n������       D                        ��������                            ���������  H@    	                        ^������`  �  �  B�  �     �             ���`���  B  �� !     �   @            ����/���   �0     � �� �            �������  1�� P     �               ��O����  ����    0 �       �    /��< <��  > <    � ?��        ?     [��� ����� $@� �ǐ      `        ~     ��� � ����( 	� �� 
 @�  �  �      �     ��� � 7���A �� t A   �       �     m�� �� �� � G �� 9 $�  8 ���       ��     _����� � ������ x���      ���    �����?����@ @ �����     ���    ��H?�����HH?���   �?��� �    ?���    ��?���/����?���0  0������    ?���    o�P��������������   1�����`    ����   ��?�z�����?�z���   s�w��p    ?$r�  ��0���K�� �����L  w�p�8    0p�  ��0� �+�� ������h   �p�    0� �  ��0�� ��7��@,������6   �� ��    0�� ��  ��x�L����@,x���   ����    x�@��  �|��������X|��3�� @ ����    |�����  ��� ��
���X�����J    �  ��    �  _�  ���������0�����݀  @�� ���    �� ���  � ��� ����� ���������  @�����    ?�� ���  ���������� �������   @?�������   ?� ���  �`ߟ������� `ߟ�!���  �?�=����   �  |�� �A��~����a￀ ����  ���?���   �  >��� �A�>�>���a�? ~��  ���ߟ�π   <  �� �A�z@�/~ ��a�z�b���  ��^�_��   x  ~ � ��������_� ����P��`  z��~#�    � x @ �����7����7�`   �����!�      0 @ ������/����X/�`   ����� �         @ ���s�������`   �_�w� �     �   @ ���(�
�����"��   ����� @         @ ��X����C�"�� � ����� @         @ ��(�
�o�C�"�p � ����� �         @ �C�S��o�C���p � �_�w� �     �   @ �C��ǈ��C�	H�` � ����� �         @ ������#��` ����� �         @ �A���п�_� S��P��` �z��  �          @ �a�zs��?¿�i������  �}\_ �    x O  � �q��.���u� .��  �}�����    <    � �?��~�¿�?��  ���  ��>���p�  �>  >  � �>߁����� >߂ �熀  ��?}�~�      |  � ��������� ����c��   @ ����    � �   �'�������� ��������  @ ���     ��   ��?������3��������  @ ��     ��   �<9���~
���X�������     C���     ���   � ~������X?��� @  ���� �      ��   �� �?���@,���U    � ��      >�    ���������@.��t��V     �  �      p    �������/�� �����l        �            ���������� ������        8            ���������	�������         8            o������ǯ��������Ǡ         p             w�@�������`������  �    `         @  �� ?�����@0?���@   �    �         @  ���������  �����   �   �    �     �  ������߀ L���=�    p        @       ��� 6���  6 ���7     8        0       ���  i��� 	�/� �                   ��� ��}�@��_ � �       p            ��`> o��   > p     �� �         `   =���� 9���  �� ��      �  �      �  �   ��������  ��ƀ    p  ?       0      �����;���    o��:        �         8    {������x  � �� �    ���       ��    ���������   ���  @     �         �     ������{�  � �  �                        ���������                                   ���������                                }�������                                   �������                                   �������   @                            �������                                                                   Q Q  g�����0   �8  �                         �?���}�   @�  �                      ~�����d   �    @�                        n������       D                        ��������                            ���������  H@    	                        ^�������`  �      B�  �     �             ���������  B      !          @            ���������            �      �            ��������   �  P                       ��������  ��      �              /����?���   �0    ��               [�������� $@ ��      �              ���� �1���(  G��� 
 @� 8 �  �      �     ���������A ��<� A   `�       �     m��`��?�� � x��0 $�  �����       ��     _�������� � ���� � ���`      ���    ������o�� 	�����  @ ���      ���    ���?������H ?���v    ?���     ?���    ��?������� &?���    �����     ?���    o���������� @���̀    9�����      ����   ���?�z���� �?�z���    s�w��     ?$r�   ��0���_�� 8����`   ��p�    0p�   ��0� ���� 0������   ��p��    0� ��  ����� ����@������p   �� ���    p�� ��@  ��x�L����@����   ����`    x�@��   �|���������	���3�� @����p    |�����   �?�� �����?�����T   �  ��    ?�  _�  �?�����S���?�����T   �� ���    ?�� ��P  ���� ����� �������   �����    ?�� ���  ����������� ������   ?������    ?� ���  ��ߟ������� ߟ�!���   ?�=���    �  |��  ����~���� -￀ ���   ��?��    �  >��  ���>�>��� -�? ~�   ��ߟ��    <  �  ���z@�/~�� -�z�b��   �^�_�    x  ~  ���������� [���P��    z��~&     � x  �����7��� [�7�     �����&       0  ������/��� [�X/�     �����&           ���s���� [���     �_�w�&      �    ���(�
��� [�"�     �����&           ���X���� [�"�     �����           ���(�
��� [�"�     �����           ���S��� [���    �_�w�      �    ����ǈ��� [�	H�     �����           �������� [��    ����           �����п��� [��P��    z��             ���zs��?��� -�������   }\_      x O   ����.��� )� .�   }����     <     ����~���� /��  ��   �>���p   �>  >   ��߁����� ߂ ��   �?}�~       |   ���������� ���c��    ���     � �   ���������� ������    ���     ��   ��?����S����������    ��8     ��   �<9���~_����������    C���0     ���   � ~���������� @ ���� �      ��   ����?�?��@����0    � ��      >�     ��������O��@���t��P     �  �      p  @  ��o������� o�����`   �   �          @  ��7�������� 7������   �    �          �  �����������������    `         @       o�)�������� �����ۀ    p                 w�����6���� V�����    8               ���?���m���@ +?���n                    ����������  �����       p            ���g���7�߀ 
g���8     �  �             ��������  �����     � �     �   �   ���FO1?��� G��q@     �0 �      @      ��y���}�@� ��΀ �    >  ?       8      ���?�1���    ~?�2       ��         0    =��������   ��       ���       ��    ��������   ��`      ?��        �     ��������     ?��                          {�������x  �      �                       ���������         @                       ������{�  �     �                        ���������                                   ���������                                }�������                                   �������                                   �������   @                            �������                                                                   Q Q  g�����0   �8  �                         �?���}�   @�  �                      ~�����d   �    @�                        n������       D                        ��������                            ���������  H@    	                        ^�������`  �      B�  �     �             ���������  B      !          @            ���������            �      �            ���������       P                       ���������                            /���������                              [��������� $@  �                         �����?����(  ��  
 @�  �   �            �����o����A  �p  A    �?�              m��������� �  8���  $�    �p         �     _��g������ �  ����  �  �        �     ��������� �����  @   ���        ���    ���3������H ?���@     ����     ���    ��O�������� ����    ����@     ���    o����������� �����     ?���       ?���    ���?�zo��� ��z��     w�      ?$r    ���������  ����    �p�      p�   ���� ����  &�����     �p�      � �   ����� �����@ L�����     ;�� ��     �� ��   ����L�����@ H���     ?����     �@��   ����������� ���3��� @ ����     �����   ��� �����������    ��  ��    �  _��  �_���������_������    ��� ���    �� ���  ����� ����  ������@   ?�����    ?�� ��@  ����������� ������   ?������    ?� ���  ��������_�� ߟ�!��@   ?�=���    �  |�@  ����~�/�� ￀ ���   ��?�`    �  >�   ��w>�>��� �? ~�   ��ߟ��    <  �  ��yz@�/~��� �z�b���   �^�_p    x  ~   ��������� ���P��   z��~0     � x  �����7��� �7�    �����0       0  ������/��� �X/�    �����0           ���s���� ���    �_�w�0      �    ���(�
��� �"�    �����0           ���X���� �"�    �����8           ���(�
��� �"�    �����8           ���S���� ���    �_�w�0      �    ����ǈ��� �	H�    �����0           �������� ��   ����0           ��~��п��� ��P��   z�� 0            ��|zs��?��� �������   }\_ p     x O    ����.?�� � .�   �}����`    �<      ����~�?�� ��  ��   |>���p`    `>  >    ���߁���_�� �߂ ��@   x?}�~�       |@  ���������� ���c��`    ����     � �@  ���������  �����@    ����     ��@  �?��������������    ����     ���  �|9���~����������    �C����     ����  ��~������� ����� @ @����       ��   ��X�?�
���@ ����z�    # � �       >�    �����������@ O��t��     0 �        p    �����������  '�����                     �����������  ;�����                    ����������� �����         0            o��?���?���� ���0     �   �             w��������� ?���`    � �         @   �����������@ �����      � �      �  �   ����������   ����     x              �������߀  x���        |            ����?�w����   ?�t       ��         p    ����������  ��      ���        ��    ��������}�@� ���  �     ?�         �     ���������     �                           =���������                                 ���������                               ���������                                  {�������x  �      �                       ���������         @                       ������{�  �     �                        ���������                                   ���������                                }�������                                   �������                                   �������   @                            �������                                                                   Q Q  g�����0   �8  �                         �?���}�   @�  �                      ~�����d   �    @�                        n������       D                        ��������                            ���������  H@    	                        ^�������`  �      B�  �     �             ���������  B      !          @            ���������            �      �            ���������       P                       ���������                            /���������                              [��������� $@                             �����������(        
 @�       �            �����������A        A                     m�������� �   �   $�                      _������� �   p�  �   �                ���� o���   p   @   ���               ����������H  ��      �`            �����������  ���      ���       ���    o�����������  o���       ���       ���    ����z�����  ��z��      ow�{       $rx    ���?w����  ?���@     �p|�      p|    ��� ����  ����     �p~@      ? ~    ���� �_���@ ���P     �� ��      � �    ����L?����@ �f�?�     ���P      �@?    ����������� 	��3��  @ ����     �����   ���� ������ �����     �  �     �  o�   ����������� �����     �� ��     �� ��   ���� �����  '����     ����     � ��   �����������  G����     ?�����     ߀ ��   ��׿�������  W��!��     /�=��     �  |�   �����~���  /�� ���    W��?�     �  >�   ��'>�>}���  �? ~}�    _��ߟ�     <  y   ���z@�/}��  �z�b��     W�^�_{�    x  y   �������?��  ���P�@    Qz��{�     � y   ��_��6��� _6�    �������       0�  ��_���.��� _X.�    ������         �  ��_s���� _��    ��_�w�      �  �  ��_(�
��� _"�    ������         �  ��X���� "~�    �������         �  ��(�
��� "~�    �������         �  ��S���� �~�    ��_�w��      �  �  ���ǈ��� 	H~�    �������         �  ��~����� ~~�    ����         �  �����н?��  ��P�@    Az���            ���zs��=��  ������     C}\_�     x O   ��1��.���  �� .�    N}����      <     �����~���  +�  ��    T>���s      >  >   ���߁������  W߂ ��     (?}�~        |
   �����������  _��c��      ���      � �   ����������  /����     ���      ��   ��?�������� /�����     ��      ��   ��9���o���� �����     C���      ���   ��~���s���� ���  @ ����       ��   ���?�����@ ����      � 0       >�    �����������@ ��t��      � `      p     ���?������  ?���`     � �         @   �����������  �����     �  �      �   �   �����������  �����      x         `      o�����������  S���       <               w���{������  <{�      � �             �����k����@  �l       ��         `    ����������   ��      ���        ��    ����O���߀   ���        ?�         �     �����������    �                           �����������                               ��������}�@�       �                       ���������                                  =���������                                 ���������                               ���������                                  {�������x  �      �                       ���������         @                       ������{�  �     �                        ���������                                   ���������                                }�������                                   �������                                   �������   @                            �������                                                                   Q Q    <�       � �       @                  �đ�      ;n        �                 >�>`      �� ��      @                  �����               @                ;��f     �l�      �                 L�?�_�     3��f      � @�               �������    @       �  �              g�����`    �   �     @                  ����?�   �   �`                        ;�����h   �    �                       �������                @              =�������                               [�������   $  ?�    @                  ��`?�v�  H��� �      �                n���o��@  � �p D�  @  ��        `     }�������`  � ���  �  ! �p B      �     ��'�p�� D ���� @   �        �     ������ @��}�     �       �     ��0���_�� <���`  � ����� �     ���    
��C�����  s��� P ����@     ���    �������� 	 �����@  ���      ���    ���z|k�� 
@��z��    w�|      $r|    +����7��  3���t    @p     p    ;�� ��� �"�����   �p�      � �   W��� ���� (�L�����   9�� ��     �� ��   W�H�L��� ( ����@  ;����     �@��   ����������	 ���3��  @ ����    �����   ���� ����B������  ��  ��    �  _�  �������?߀P�����    ��� ���    ?�� ��   ����� ��_� R������` ��?�����    �� ��@  {�������_��������@  ?������    � ��@  _�������ߟ�!��  �=���    �  |�   [����~�/������ ��0   ��?��    �  >�   ��7>�>~�� �? ~~�����ߟ�p    <  ~   ��9z@�/~��@�z�b��� �^�_~p    x  ~   ��?�������H���P��   z��~0     � x  ����7W��H7X    �����0       0  �����/_�� X/X	 H �����0           ��s�_��H�X    �_�w�0      �    ��(�
_��H"X    �����0           ��X�_�� "X	 H �����0           ��(�
_��H"X    �����0           ��S�_��H�X    �_�w�0      �    ���ǈ_�� 	HX	 H �����0           ��~��_��H~X   ����0           ��>��о���H��P��   z�� 0            ��<zs��>��@������� }\_ p     x O    ��!��.�� !� .����}����p     <      [���~�������  ��   |>���p`    `>  >    _��߁���O�߂ ��P 8?}�~�       | @  {�������������c��`   ����     � � @  �������_� R �����` �� ����     �� @  ��?�����߀P������   ����     �� �  ��|9���~���B������  �C����     ��� �  ���~������	 ����� @ @����       ��   W�X�?��� ( ����z @  # � �       >�    W�������� (�]��t��     �        p    ;������� �&�����                    +��?���o�� @���l                    ��������� 
 �����         0            ��G������  O����     �   `             ���������  �����   @  @         @   ������x  ������ �    � �      �  �   ����r���   ��r�     x               ����ǎ���   X��       ? |             ����u���  ! 7�v B     ��         p    ��������  @ ��      ���        ��     ���������    ���        �         �      w�������   @ �                          /�������                                �������         @                         �������                                  �������                                   �������     @                             w�����@    �  �                          ~���      � @�                           /��o��      �                            �����       @                           �����      @                              ��o��       �                             ;���       @                                                          Q Q    <�       � �       @                  �đ�      ;n        �                 >�>`      �� ��      @                  �����               @                ;��f     �l�      �                 L�?�_�     3��f      � @�               �������    @       �  �              g�����`    �   �     @                  ����?�   �   �`                        ;�����h   �    �                       �������                @              =�������                               [�������   $        @                  ������v�  H�     �                        n������@  �  �  D�  @                   }��0��`  �  ��  �  !  �  B             ����o�� D �p @    ���        �     �������� @ ��     �`       �     ���������  3���   � ���  �    ���    
��O�����   ���� P  7���      ���    ��������� 	 �����@   ���      ���    ���z}_�� 
@�z�`     �w�~�      ?$r|    +��������  �����    @p`     p    ;�� ��� ������   �p�      � �   W��� ���� (������   �� ��     �� ��   W���L���� ( 2��� @  ����     �@��   ����������	 $�3��  @ ����     ~����   ���}� �����B D}����   ?�  �     }  _�   ���?�����߀P N?����    ?�� ��     ?� ��   ��O?� ���� R �?����  �� ?����     ?� ��   {����������� ������   _�����     � ��   _������� ���!��   _�=���    �  |�   [�o��~����o�� ��@    ���?��    �  >�   ��w>�>�� w? ~��� ���ߟ��    <  �  ��yz@�/~��@yz�b���  ��^�_�    x  ~�  ���������H��P��    �z���     � x�  �����7_��H�7`    ������       0@  ������/�� �X/`	 H ������         @  ���s���H��`    �_�w��      �  @  ���(�
��H�"`    ������         @  ���X�_�� �"@	 H ������         @  ���(�
_��H�"@    ������         @  ���S���H��`    �_�w��      �  @  ����ǈ�� �	H`	 H ������         @  �������H �@   �����         @  ��~��о���H~�P��    �z���          �  ��|zs��>��@|������  �}\_�     x O �  ��a��.��  a� .��� �}����    @<   �  [�c��~����� c�  ��    �>���q�     >  > �  _��߁��� �߂ ��   X?}�~�       |   {�?�������� ���c��   @���      � �   ��������� R _����  ��  ���      ��   ���?�����߀P _�����     ��      ��   ���9���u���B /�����   C���      ���   ���~������	 /���  @ ����       ��   W���?��� ( ���h @   � �       >�    W�������� (���t��    � 8      p    ;�������� �
�����      p             +�����O�� @���P    �   �         @   ��������� 
 �����     �  �      �   �   ��O���?��  O���@      �  �      @      ��3�����   ����    |        0      ������x  � ,���  �     |             ����g���   �h      ��         `    ���t���   t        ���        p     ���������  !  O�  B      ?�         �     ���������  @  �                           ���������                                   w�������   @                             /�������                                �������         @                         �������                                  �������                                   �������     @                             w�����@    �  �                          ~���      � @�                           /��o��      �                            �����       @                           �����      @                              ��o��       �                             ;���       @                                                          Q Q    <�       � �       @                  �đ�      ;n        �                 >�>`      �� ��      @                  �����               @                ;��f     �l�      �                 L�?�_�     3��f      � @�               �������    @       �  �              g�����`    �   �     @                  ����?�   �   �`                        ;�����h   �    �                       �������                @              =�������                               [�������   $        @                  ������v�  H�     �                        n�������@  �      D�  @                   }�������`  �       �  !      B             �������� D      @                      ���0��� @  ��      �               ����_���  �`   �  ���  �     �     
���������   ���  P  �`       �     ��������� 	  3��� @   �       �     ����zr��� 
@ o�z�      w�l       $r`    +��_��}��   �����    @ 'pr      pp    ;�? ~?�� �?���@    �p}�       |    W�� ��� (����    �� ��      ?� �    W����L���� ( ���� @  ��`      �@�    �����������	 ��3��  @ ����      �����   ���}� �����B }����   �  �     }  _�   ��������߀P ����    �� ��     � ��   ��� ���� R �����  �� ����     �� ��   {����������� '����    �����     � ��   _����� /��!��   �=��     �  |�   [����~����� _�� ��     '��?�     �  >�   ���>�>~��  W? ~ �� /��ߟ�     <  ~   ���z@�/��@ Yz�b��   '�^�_~     x  ~   ��߄������H _��P�     !z��      � ~   ��?��7��H �7�    @�����        3   ��?���-��  �X-�	 H @�����         !   ���s����H ���    @�_�w�       �    ���(�
���H �"�    @�����            ���X����  �"}�	 H @�����            ���(�
���H �"}�    @�����            ���S����H ��}�    @�_�w�       �    ��?�ǈ��  �	H}�	 H @�����            ��>����H �}�    A����            ��^��к��H ޅP��    !z��             ���zs��;��@ \�����   #}\_      x O   �����.��  Q� . �� .}����      <     [����~����� [�  �     $>���~      >  >   _��߁���� /߂ ��   ?}�~        |   {����������� /��c��    ���      � �   ��������� R ����  �� ���      ��   ���?�����߀P �����    ��8     ��   ���9���S���B �����   C���8     ���   ���~���/���	 ���  @ ����p      ��    W��?�W�� ( ��X @  �� �      >� @   W�?���o�� (�?�t�p   ���      p @   ;�������� ������    � �      �  �   +�������� @�����     x                ��S����� 
  ����      <               ���{����   l�       � �             ����k���   �l     ��         `    ������x  � ��  �    ���        ��    ���������   ���       ?�         �     ���������    ?�                           ���������  !      B                        ���������  @                               ���������                                   w�������   @                             /�������                                �������         @                         �������                                  �������                                   �������     @                             w�����@    �  �                          ~���      � @�                           /��o��      �                            �����       @                           �����      @                              ��o��       �                             ;���       @                                                          Q Q    <�       � �       @                  �đ�      ;n        �                 >�>`      �� ��      @                  �����               @                ;��f     �l�      �                 L�?�_�     3��f      � @�               �������    @       �  �              g�����`    �   �     @                  ����?�   �   �`                        ;�����h   �    �                       �������                @              =�������                               [�������   $        @                  ������v�  H�     �                        n�������@  �      D�  @                   }�������`  �       �  !      B             �������� D      @                      ��������� @                            ��������   �    �       �            
��������    p   P   �               ��������� 	  ��� @                     ����z/��� 
@ �z�      w�@        $r     +��������   ���     @ pp       p     ;�� u��� � 3���     pH        @    W��� ���� (� G���     ?� �       � �    W���L��� (  ���� @   ��       �@�    ������?���	 �3�@  @  ����      ���    ���=� ߟ���B =��ߠ    �  ~�      =  ^�   ������_�߀P ���@    �� ��      � �@   ����� ���� R �����  �� ����      �� ��   {����������� ����    �����      � ��   _������ 	��!��   �=��     �  |�   [����~����� 	�� ��     ��?�     �  >�   ���>�>o��  ? ~h �� ��ߟ�     <  h   ���z@�/o��@ z�b��   �^�_x     x  h   ����������H ��P�     	z��|      � h   �����7���H 4     �����        4   ������%���  /X& 	 H �����         $   ���s����H /�     �_�w�       �    ���(�
���H /"     �����            ���X����  /"v 	 H �����            ���(�
���H /"v     �����            ���S����H /�v     �_�w�       �    ����ǈ���  '	Hv 	 H �����            ��������H (v     ����            �����Ы���H �P�     z��             ���zs��+��@ �����   }\_      x O   ����.��  � . �� }����      <     [����~����� �  �     >���x      >  >   _��߁���� ߂ ��   ?}�~0        |   {����������� ��c��    ���p      � �    ��������� R ����  �� ���`      ��    ���?���_�߀P ���@    ����      ��@   ���9��؟���B =��ޠ    �����      ����   �����������	 ����  @  �����      ����   W��O?�y�� (  Ͼ�y� @   p�       @>�    W�������� (� w�t�     8�       0p    ;�������� � )���      <             +���w�3��� @ w�4      � �         0    ��������� 
  ���       ��       � �    ���p?���   p@        ���        p     ���������    O�       ?�         �     �������x  �  �   �                       ���������                                ���������                                 ���������  !      B                        ���������  @                               ���������                                   w�������   @                             /�������                                �������         @                         �������                                  �������                                   �������     @                             w�����@    �  �                          ~���      � @�                           /��o��      �                            �����       @                           �����      @                              ��o��       �                             ;���       @                                                          