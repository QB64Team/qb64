�l  �z��                 `                                              `                                              `                                              `                                             �` 0                                           �` 0                                           �` 0                                           �` 0                                            ` 0                                            ` 0                                            ` 0                                            ` 0                                           g�8<��ny����<��<                               g�8<��ny����<��<                               g�8<��ny����<��<                               g�8<��ny����<��<                               3lٰf��l��m���f                               3lٰf��l��m���f                               3lٰf��l��m���f                               3lٰf��l��m���f                               �o�0f�������0>͛~                               �o�0f�������0>͛~                               �o�0f�������0>͛~                               �o�0f�������0>͛~                                                                                                                                       �l03f�����͛0f͛`                                                                                                                                                                                           �lٰ3f́�l͛m�0f͛f                                                                                                                                                                                           g�<���fy���0>��<�                                                                                                                                                                                                                                                                                                                                                                                                                           �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ?��                ��                ��                                                                                                                                                                       � |                �               | �                                                                                                                                                                      x  �             �                �  <                                                                                                                                                                     �   8                 �             8   �                                                                                                                                                                                     0                 �    `                                                                                                                                                                    0    �            �                                                                                                                                                                                         �     `                �                                                                                                                                                                                                          `           0     �                                                                                                                                                                                   0                 �      `                                                                                                                                                                                   @                                                                                                                                                                                                 �          �                                                                                                                                                                                         �       `                �                                                                                                                                                                                                          @                                                                                                                                                                                                                             �                                                                                                                                                                                                  @        @                                                                                                                                                                                                   �                                                                                                                                                                                          @                                                                                                                                                                                                   �        �                                                                                                                                                                                         @         @                                                                                                                                                                                                 �                           �                                                                                                                                                                                                         @                                                                                                                                                                                                                           �                                                                                                                                                                                                          �                                                                                                                                                                                              @          @                                                                                                                                                                                              �                                                                                                                                                                                      @                                                                                                                                                                                                      @                                                                                                                                                                                                 �      �                                                                                                                                                                                                �      �                                                                                                                                                                                    @           @                                                                                                                                                                                       @     @           @                                                                                                                                     @                                                   �     �                             �                                                                                                                    �            @                  @                        �                             �                                                                             @                  @                               @                  �                                                    @                                                                             @                  �                               �                  �                                                    @                                                                             �                  �                               �                                                                                         �                                                            �                                                                                                                                          �                                                                                                                                                                                                       �                                                                                                                                                  @                                       @            @                                                                                                @                                                 �                                       @            @                                                                                                �                                                                                        @            @                                                                                                                                                                                        @            @                                                                                                                                                                                          �                                                                                                                                                                                                       �                                                                                                                         �                 �                 �                                        �                    �                  �                                                                                �                 �                              `                           �      �                              �                                                                                  �                 �                              @                           �     �                             	�                                                                                  <                 �                 p            �          @                     �                            �                 0                                                                                 �                 �            �          @                                 4                 �                 `                                                                s�                7�                 1�           �          @                                 #                 '�                  �                                                                ��                /��                c�                     @                    0           l�                3                 A�                                                                �<                _��                ���           �         @                     8           _0                N|�                �s                                                                ��                ��<               ���           0         @       �              p           ��                �0               ��                                                               ���               ���               �<                    @     @ 0              � �          ��                <��               �0                                                               ���              ���              ?��                    @     �              � 0          ���              9��               ��                                                               3��<              ���              ���           �        @     �              �           !�0              y���              7��                                                               7���              ���<              ����           0        @       �                        #��               ���0              o���                                                              g����             ��?�              1���<                   @       0               �         B���              ��?�               ���0                                                              ����             ����             #��?�                   @                      0         �<��             	���              ��?�                                                              �� �<             ����             ߀��        0   �       @                               �� �0             ����             ��                                                              �� ?�             �� �<             ���        !   0       @       �                       �� ?�             �� �0             ����                                                            x ��            �� ?�             '�� �<        `�         @        0               �        	x �             �� ?�             ׀ �0                                                             ?x ��            �� ��            @�� ?�         �                         �        0         x ��            5� �              ׀ ?�                                             @              #�  �<            N� ��            �;� ��        @   �                      �                 �  �0             J� ��             +� �                                             �              A�  ?�            �  �<            � ��        @   0                �      �                  �  ?�             �  �0             � ��        @                                                 @�  ��           x  ?�            �  �<                         �   0      �         �         ^  �             x  ?�             �  �0        @                                                 ��  ��            x  ��           �  ?�                         �         �         0         ^  ��            x  �             �  ?�        �                                                  �o   �<            �  ��           �  ��           �           @         @          @       /   �0             �  ��            �  �        �                                                  o   ?�           @�   �<           �  ��           0           @    �     @          @       /   ?�             �   �0            �  ��                        @                                7�  ��          � �   ?�            x   �<                           0     @      �    �@       �  �             ^   ?�            x   �0                        �                                 7�  ��          � �   ��         @ x   ?�                                @      �    0@       �  ��            ^   �            x   ?�                        �                 @               �����0           o������         � ������            �                            @    �       �  ��0            /  ���            �  ��                                         �               ������           o�����           ������            8                �            @    �       ������            /�����             ������                                                           ��           4   ��           �  ��       ����            ����              /���  �          ��               ��            P  ��                                                        ������           7������           ������                            @                        ������            ������            _�����                                                        ������           ������           o�����                            @                       ������            ������            /�����                                                        ������           �����            o�����  �                           �                       ������            �����             /�����                                                        �����           �����             7�����  �      �                     �                       �����            �����             �����                                                          x                 �             @   7�      @      �    @                                       x                 �                 �                                              @                 �                 �             �   �      @      @    @                                        �                 �                 �                                              �               @ �              @  �                �             @    �      �                                  �                 �                 �          @                 @                                @  �              �  x                �                  �      �      �                            ^                 x                 �          @                 �                                �  �              �  x                �                       @      �                            ^                 x                 �          �                 �                                �  o                �                �                      @      @                            /                  �                 �          �                                                   o                �                �                             @          �                   /                  �                 �                                                             7�                �                 x                                       @      �   @         �                 ^                 x                                                              7�                �            @    x                                               �   �         �                 ^                 x                                           @                  �                o            �    �                                              @   �         �                 /                  �                                           �                  �                o                �                               @             @            �                 /                  �                                                             �                7�                �       �                         �                          �                 �                 ^                                                             �                 7�                 �       @        @                                          �                 �                 ^                                                               �                 �                 o                �        �                                 �                 �                 /                                                               �            @    �                 o                       @                                 �                 �                 /                          @                                    x            �    �                 7�            �                           �                  x                 �                 �                         �                                     x            �    �                 7�            �                          @       @          x                 �                 �                          �                                     �                �                 �            @                                   �           �                 �                 �                                                           @   �                �                 �            @                 @                           �                 �                 �        @                                                  @    �                 x                 �       �       `               ��                           ^                 x                 �        @                                                   �    �                 x                 �               �          �     �                            ^                 x                 �        �                                                   �    o                 �                 �                       @     @                            /                  �                 �        �                                                       o                 �                 �                       0     @           �     `            /                  �                 �                                                                7�                 �                 x                             `           0     ��            �                 ^                 x                                                                 7�                 �                 x        �    `                !�                �             �                 ^                 x                                                                                   h                 �        0    �            �                     X             
                  (                  �                                                                                   `                 �                         0                 �    `                                                  �                                                                                                                �   8                 �             8   �                                                                                                                                                                     x  �             �                �  <                                                                                                                                                                      � |                �               | �                                                                                                                                                                       ?��                ��                ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      � `�  ��         ̀`             �         0                                                                                                                                                              0    ��         l `�             0     0                                                                                                                                                                 0    ��          `�             0     0                                                                                                                                                                 1�n�><��;`<��<     �|�y�<��y�      ��͹��3π                                                                                                                                                            1��lٻ�����f     ͳv�Ͷf���      ͳ3m�m�7m�n�                                                                                                                                                            1��lٳ>����>͛~      m�f���~��͘      3?m��3�f6l�                                                                                                                                                            1��lٳf����f͛`      m�f���`�f͘      30m�3c6l�                                                                                                                                                            1��lٳf���`f͛f     m�f�ͶfͶ͘      �3m�m�6m�l�                                                                                                                                                            1��f�3>��30>��<     ͟f`y�<��y�      �m�͙�g3��                                                                                                                                                                                                                                                                                                                                                                                      �        >                                                                                 