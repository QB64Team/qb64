��g  �-            �6  00�  �                         �6  00�  �                         �6  00�  �                         �6  00�  �                         �6  0x   �                         �6  0x   �                         �6  0x   �                         �6  0x   �                         ff  0x   �                         ff  0x   �                         ff  0x   �                         ff  0x   �                         fgǏ00>>y���>                       fgǏ00>>y���>                       fgǏ00>>y���>                       fgǏ00>>y���>                       fglٰ0��f́���                       fglٰ0��f́���                       fglٰ0��f́���                       fglٰ0��f́���            �����������               ����������������������               �����������           ?�o߰~�f�����                                                                                                                                         ?�l0l3f����3                                                                                                                                         �lٰl�f́���                                                                                                                                         �g�0>3>y���>                                                                                                                                                       0                                                                                                                                                       0                                                  