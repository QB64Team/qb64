�&^  �k 6              ��������������              �              ��������������                          �              ��������������                          �              ��������������                          �              ��������������                          �              ��������������                          �              ��������������                          �              ��������������                          �              ��������������                          �              ��������������                          �              ��������������                          �              ��������������                          �              ��������������    @                    �              ��������������                       �              ��������������                       �              ��������������X͢sNX�                  �              ��������������e)"�Qe                   �              ��������������D�"�QD�                  �              ��������������DI"�QD@                  �              ��������������E)&�QE                   �              ��������������D�qND�                  �              ��������������                          �              ��������������                          �              ��������������                          �              ��������������                          �              ��������������                          �              ��������������                          �              ��������������                          �              �������������� !   y                    �              �������������� !  @�                    �              �������������� Q  @�                    �              �������������� Q�`�c�x�                �              �������������� �Q@��QE                �              �������������� �Q@�QE�                �              �������������� �Q@�QE                �              ��������������S@�QE                �              ��������������� y�x�                �              ��������������       @                 �              ��������������       @                 �              ��������������                          �              ��������������                          �              ��������������                          �              ��������������                          �              ��������������                          �              ��������������                          �              ��������������                          �              ��������������                          �              ��������������                          �              ��������������                          �              ��������������                          �              ��������������                          �              ��������������              ��������������              �������������              �������������              �������������              �������������              