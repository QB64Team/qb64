��]  T4]                                    ������������������������������������                                    �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������        ~`         �                        ~`         �              �         ~`         �               ������������������������������������        c`     `  �                        c`     `  �              �         c`     `  �               ������������������������������������        c`     `  �                        c`     `  �              �         c`     `  �               ������������������������������������        cg�x>s���<�?�                   cg�x>s���<�?�         �         cg�x>s���<�?�          ������������������������������������        ~l����fl ��f��ـ                  ~l����fl ��f��ـ        �         ~l����fl ��f��ـ         ������������������������������������        `oϘ��g���~϶߀                  `oϘ��g���~϶߀        �         `oϘ��g���~϶߀         �����������s?�̙��>d��&I'�����������                                            `l��3f��`ٶ�         �                                    ����������&I3�L���>d��&I&����������                                            `lٶ��fl��fٶـ        �                                    ����������pc����3�>d��0I0�����������                                            `g��x33���<϶�         �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������� �_��������������                                     }       0߀��   �     ���  �                                    ������������O'?�_����������������                                             ��� ��   �    �@  �                                    ������������F'?�_����������������                                             ��� ��   �    �@  �                                    ���Li͍?�F'=�_?�c��t�'c�m�����                                     c�䳖2r����J���q�x�9��r�@  �                                    ���k��[��t��� }�_u���]w�u���]�m�����                                     �A�YJ� ?߂J�� 
(���E$�
�@  �                                    ����>�.�u��@'�U_t��Aw�u��_�m�����                                     ��'�"� ������z(���E$��z�@  �                                    ���������u��I'�U_u�u�_w�u���_um�����                                     $� ����� �(��"�E%���@  �                                    �����[��u��I'��_u�u�]w�e���]us�����                                     A�QJ� ���� �(��"�E%���@  �                                    ����ln͍� �'��_?�c����c�w�����                                     �䓑2r �0����y�xi9$�z�@  �                                    ������������������������������������                                                                 @  �                                    �����������������������������������                                                                 0�  �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                        ?����������������������      �                                    ������������������������������������                                                                     �                                    ������������������������������������                                                                     �                                    ������������������������������������                                                                     �                                    ������������������������������������                                                                     �                                    ������������������������������������                           A              ����������������������      �                                    ������������������������������������      ���������������������              ����������������������      �       ���������������������       ������������������������������������      ���������������������              ����������������������      �       ���������������������       ������������������������������������      ���������������������              ����������������������      �       ���������������������       ������������������������������������      ���������������������              ����������������������      �       ���������������������       ������������������������������������      ���������������������              ����������������������      �       ���������������������       ������������������������������������      ���������������������              ����������������������      �       ���������������������       ������������������������������������      ���������������������              ����������������������      �       ���������������������       ������������������������������������      ���������������������              ����������������������      �       ���������������������       ������������������������������������      ���������������������              ����������������������      �       ���������������������       ������������������������������������      ���������������������              ����������������������      �       ���������������������       ������������������������������������      ���������������������              ����������������������      �       ���������������������       ������������������������������������      ���������������������              ����������������������      �       ���������������������       ������������������������������������      ���������������������              ����������������������      �       ���������������������       ������������������������������������      ���������������������              ����������������������      �       ���������������������       ������������������������������������      ���������������������              ����������������������      �       ���������������������       ������                     >��������      ����������������������                                          �                                    ������������������������������������                                                                     �                                    ������������������������������������                                                                     �                                    ������������������������������������                                                                     �                                    ������������������������������������                                                                     �                                    ������                      ��������     ?����������������������                                          �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                                                      �                                    ������������������������������������                                    ������������������������������������                                    ?�����������������������������������                                    ?�����������������������������������                                    ?�����������������������������������                                    ?�����������������������������������                                    