��_  ܽX�                                                                            ���������������������������������������������������������������������������                                                                                                                                                      ���������������������������������������������������������������������������                                                                                                                                                                                                                                 ���������������������������������������������������������������������������                                                                                                                                                                                                                                 ���������������������������������������������������������������������������                                                                                                                                                    �                                                                           ���������������������������������������������������������������������������                                                                         ��                                                                                                                                                  ��������������������������������������������������������������������������
�                                                                       P@                                                                       �                                                                           ������������������������������� ��������?����������������������������������                                                                       �@                             ��       �                               H                                                                           ���������������������������������?����<����������������������������������                                                                       p@                             �� �   ?À                               �                                                                           �������������������������������O�������8���������������������������������                                                                         ��                            �x �  ;ǀ                                                                                                          ����������������������������������������8���������������������������������                                                                                                        <    qǀ                                �                                                                           �������������������������������������������?������������������������������                                                                                                         <     q�   �                                                                                                         ��������������������������������������������������������������������������                                                                                                         8<   < x  �                                                                                                         ������������������������������������� ?����8?������������������������������                                                                                                         x?��8��                                                                                                         ����������������������������������������0?������������������������������                                                                                                         p9�<�� <<��                                                                                                         �������������������������������0������8������������������������������                                                                                                         ���=�� �y��                                                                                                         �������������������������������<p�����0������������������������������                                                                                                          �Ï?�� ����                                                                                                         ������������������������������� �`����0������������������������������                                                                                                          ��~�� ����                                                                                                         ���                           ���������������                          ��  ����������������������������� �8<�� x�x?���������������������������                                                                                                                                                        ���������������������������������������������������������������������������                             ��8�� y�p                               ����������������������������              ���������������������������                                                                             ���������������������������������������������������������������������������                             �<1�� <y�p                                                                                                                                                                                   ���������������������������������������������������������������������������                             �8q���8y��                                                                                                                                                                                   ���������������������������������������������������������������������������                             ��p����x0��                                                                                                                                                                                   ���������������������������������������������������������������������������                             ��` ��  00                                                                                                                                                                                     ���������������������������������������������������������������������������                             �    �     <                                                                                                                                                                                    ���������������������������������������������������������������������������                             �           <                                                                                                                                                                                    ���������������������������������������������������������������������������                                                                                                                                                                                                                              ���������������������������������������������������������������������������                                                                                                                                                                                                                              ���������������������������������������������������������������������������                                                                                                                                                                                                                              ���������������������������������������������������������������������������                                                                                                                                                                                                                               ���������������������������������������������������������������������������                                                                                                                                                                                                                               ���������������������������������������������������������������������������                                                                                                                                                                                                                               ���������������������������������������������������������������������������                                                                                                                                                                                                                               ���������������������������������������������������������������������������                                                                                                                                                                                                                               ���������������������������������������������������������������������������                                                                                                                                                                                                                               ���������������������������������������������������������������������������          �                       �    �   0     �                        �                       �    �   0     �                         �                       �    �   0     �              ���������������������������������������������������������������������������          6                       0       0   �  �                        6                       0       0   �  �                         6                       0       0   �  �              ���������������������������������������������������������������������������                                         0   �  �                                                       0   �  �                                                        0   �  �              ���������������������������������������������������������������������������          ǟ<�c�x�<�              ���g��fp;�����<y�s�                      ǟ<�c�x�<�              ���g��fp;�����<y�s�                       ǟ<�c�x�<�              ���g��fp;�����<y�s�            ���������������������������������������������������������������������������          `ݳf��`͛f�              �m�6`ٳf�36�6��6�fͳf�                      `ݳf��`͛f�              �m�6`ٳf�36�6��6�fͳf�                       `ݳf��`͛f�              �m�6`ٳf�36�6��6�fͳf�            �����     ���������������    ��      ?������������������������     �����    ������gٳ~ۇ���f�?����� �������7���ٳf`36����`ͳc ������               gٳ~ۇ���f�               7���ٳf`36����`ͳc                        gٳ~ۇ���f�               7���ٳf`36����`ͳc             �������������&L��$9�>d�?�����������������|��3&L����'�9$�s�2L�������������    �                                                                      �����lٳ`�� ��f������ �������6��ٳf036����`ͳa��������                                                                                �����������ɓ&L��$��2d�?���������������ɒd��s&L�'��'�<d�'�2L�?������������    �                                                                            6lٳf�f`͛f�              6m�6�ٳn�36�6Û6�fͳf�                                                                                       ������������&`��d�?��?���������������3�x&a����'��gÆa�������������    �                                                                            �gٟ<�3�x�<�              �����ٞ>p6�c�<y�c�                                                                                       ��������������������������������������������������������������������������    �                                                                                                                                                                                                                     ��������������������������������������������������������������������������    �                                                                                >                                                                                                                                     ��������������������������������������������������������������������������    �                                                                                                                                                                                                                       ��������������������������������������������������������������������������    �                                                                                                                                                                                                                       ��������������������������������������������������������������������������    �                                                                                                                                                                                                                       ��������������������������������������������������������������������������    �                                                                                                                                                                                                                       ��������������������������������������������������������������������������    �                                                                                                                                                                                                                       ��������������������������������������������������������������������������    �                                                                                                                                                                                                                       ��������������������������������������������������������������������������    �                                                                                                                                                                                                                       ��������������������������������������������������������������������������    �                                                                                                                                                                                                                       ��������������������������������������������������������������������������    �                                                                        ���        ����            ���           ����                                                                                                ������������������������������������������������_������������������    �               �                           �                              <�    �   �              �   �@ @  �   �    �                                                                                         �������������������������������������}������?�������������������������    �               �                           �                              "�    �   @              �     �  �        �                                                                                         �������������������������������������}��������������������������������    �               �                           �                              "�    �   @              �      @  �        �                      ��        ��             ���           ��                      ������������c����������4�������������}�N?ܢ������������c?�������������    �               �                           �                              "�r@   �   Y�p           �s��#]�@  �   ';��                     ��        ��             ���           ��                      ������������}u���������]w���������������ݭ���������[]�]]�������������    �               �                           �                              <���   �   P,��           �
J "R@@  �    �����                     ��        ��             ���           ��                      ������������a|���������]������������}��ݭ���������[A��]�������������    �               �                           �                              "��    �   Q��           �zK�"R@@  �   '��"��                     ��        ��             ���           ��                      ������������]}���������]������������}u��ݭ���������[_��]�������������    �               �                           �                              "���   �   R(��           ��J "R@@  �   (��"��                     ��        ��             ���           ��                      ������������]u����������]w������������}u��ݭ���������[]�]]�������������    �               �                           �                              "��@   �   R(��           ��J "R@@  �   (�����                     ��        ��             ���           ��                      ������������a���������na�������������}��?ݭ���������[c��c�������������    �               �                           �                              <�r    �   ��p           �zI�"R@@  �   '����                                                                                        ������������������������������������������������������������������������    �               �                           �                                     �                            �                                                                                                   �������  ���������  �������������  ������������  ���������������������    � ���        ���          ���           ���                                     �      <                      �                                                                                                   ��������������������������������������������������������������������������    �                                                                                                                                                                                                                       ��������������������������������������������������������������������������    �                                                                                                                                                                                                                       ��������������������������������������������������������������������������    �                                                                        ���        ����            ���           ����                                                                                                ��������������������������������������������������������������������    �               �                           �                                    �    (             �   �@ �  �   �                                                                                            ��������������������������������������}���������������������������������    �               �                           �                              !      �    (             �       �   @                                                                                           ��������������������������������������}���������������������������������    �               �                           �                                     �   @(             �        �                            ��        ��             ���           ��                      �����������ߘ�O�������x�6�������������}�N?ܢ���������'f3o���������    �               �                           �                               g�   �   �)�            �s��#]�  �   vy9��̐8��                ��        ��             ���           ��                      �����������ط]7��������U�����������������ݭ������������o�����������    �               �                           �                              'H��   �   �)            �
J "R@   �   IEE%P(�E                ��        ��             ���           ��                      �����������ްAw��������U�_������������}��ݭ�����������o�����������    �               �                           �                              !O��   �   �*�           �zK�"R@@  �   IE}%�Q�A                ��        ��             ���           ��                      �����������޷�w����������_������������}u��ݭ������������o�����������    �               �                           �                              !H �   �   **�           ��J "R@�  �   IEA%R(�A                ��        ��             ���           ��                      �����������ܷ]w��������Uۿ������������}u��ݭ��������������ן�����������    �               �                           �                              #H��   �   �$@           ��J "RA   �   QIEE%R(`E                ��        ��             ���           ��                      �������������w���������;�������������}��?ݭ�������q���������������    �               �                           �                              G�   �   )�@           �zI�"RA�  �   �Iy9$�I�@8��                                                                                   ������������������������������������������������������������������������    �               �                           �                                     �                             �      @     @                                                                                      �������  ���������  �������������  ������������  ��������������������    � ���        ���          ���           ���                                     �                             �      @    �                                                                                      ��������������������������������������������������������������������������    �                                                                                                                                                                                                                       ��������������������������������������������������������������������������    �                                                                                                                                                                                                                       ��������������������������������������������������������������������������    �                                                                        ���        ����            ���           ����                                                                                                ����������������������}������������������������������������������������    �               �                           �                              <�     �   �                       �   (                                                                                              ������������������������������������������������w�������������������    �               �                           �                              "�     �   ��            �         �   �                                                                                              �����������������������������������{���������������������������������    �               �                           �                              "�     �   D��            �        �                              ��        ��             ���           ��                      ������������]����������M1�������������{���������������������������������    �               �                           �                              "�p    �   D��            �        �   *'0                         ��        ��             ���           ��                      ������������]w���������5n�������������z�2P������������_�����������������    �               �                           �                              <��    �   Dʑ            �Xͯ+    �   *(�                         ��        ��             ���           ��                      ������������]��������Wu`����������������S]��������V�_�����������������    �               �                           �                              "��    �   ���            �e)(��    �    �O�                         ��        ��             ���           ��                      ������������]��������Wuo�������������~�v�W]��������V�������������������    �               �                           �                              "��    �   ���            �D�(��    �    �H                          ��        ��             ���           ��                      ������������Yw���������un�������������~���W]��������Ww_�����������������    �               �                           �                              "��    �   ��            �DI(��    �   ���                         ��        ��             ���           ��                      ������������e����������u��������������~���W]���������x������������������    �               �                           �                              <�p    �   �N            �E)(��    �   (�                                                                                             ��������������������������������������~�:��a����������������������������    �               �                           �                                     �                   �D�/(�    �                                                                                                   �������  ���������  �������������  ������������  ���������������������    � ���        ���          ���           ���                                     �                           �                                                                                                   ��������������������������������������������������������������������������    �                                                                                                             <                                                                                                        ��������������������������������������������������������������������������    �                                                                                                                                                                                                                       ��������������������������������������������������������������������������    �                                                                        ���        ����                           ����                                                                                                ����������������������������������������������������������������������    �               �                            �                               �     �     @                       �   �A                                                                                             ���������������������_�������������������������������������������������    �               �                            �                               �     �   � @                       �   @A                                                                                             �����������������������������������������������������������������������    �               �                            �                              1�     �     @                       �    A                          ��        ��                            ��                      ������������c1Ɵ�������q�����������������������������������������������    �               �                            �                              1��9`  �   3�@                       �   O                          ��        ��                            ��                      ������������}n�o������ۮ����������������������������.�������������������    �               �                            �                              *��E�  �   $Q@                       �   	�Q                          ��        ��                            ��                      ������������an��������X ������������������������������������������������    �               �                            �                              *��E  �    ��@                       �   QQ                          ��        ��                            ��                      ������������]n��������[������������������������������������������������    �               �                            �                              $��E  �    �@                       �   QQ                          ��        ��                            ��                      ������������]n��������[�����������������������������.�������������������    �               �                            �                              $��E  �   �Q@                       �   �Q                          ��        ��                            ��                      ������������aq���������q������������������������������������������������    �               �                            �                               ��9  �   �@                       �   NO                                                                                             ������������������������������������������������������������������������    �               �                            �                                     �                              �                                                                                                   �������  ���������  ����������������������������  ���������������������    � ���        ���                         ���                                     �                              �                                                                                                   ��������������������������������������������������������������������������    �                                                                                                                                                                                                                       ��������������������������������������������������������������������������    �                                                                                                                                                                                                                       ��������������������������������������������������������������������������    �                                                                        ���        ����            ���           ����                                                                                                ����������������������������������������������������}������������������    �               �                           �                              >     �   �A                       �   �                                                                                             ��������������������������������������{�������������������������������    �               �                           �                              !     �   @A             � |       �   ��                                                                                            ��������������������������������������;�������������������������������    �               �                           �                              !     �    A             �        �   D��                         ��        ��             ���           ��                      ������������������������������������;��������������M1�����������������    �               �                           �                              !8�    �   O             �        �   D��                         ��        ��             ���           ��                      ����������������������.���������������[�Q?����������5n�����������������    �               �                           �                              >E    �   	�Q             ����     �   Dʑ                         ��        ��             ���           ��                      �����������ނ�������������������������Z�������������Wu`�����������������    �               �                           �                              !}    �   QQ             �)      �   ���                         ��        ��             ���           ��                      �����������޾�������������������������j�������������Wuo�����������������    �               �                           �                              !A    �   QQ             �)      �   ���                         ��        ��             ���           ��                      �����������޺���������.���������������r��������������un�����������������    �               �                           �                              !E    �   �Q             �)      �   ��                         ��        ��             ���           ��                      �������������������������������������r��������������u������������������    �               �                           �                              !8�    �   NO             �)      �   �N                                                                                            ��������������������������������������{��������������������������������    �               �                           �                                     �                   ��)      �                                                                                                   �������  ���������  �������������  ������������  ���������������������    � ���        ���          ���           ���                                     �                             �                                                                                                   ��������������������������������������������������������������������������    �                                                                                                                                                                                                                       ��������������������������������������������������������������������������    �                                                                                                                                                                                                                       ��������������������������������������������������������������������������    �                                                                                                                                                                                                                       ��������������������������������������������������������������������������    �                                                                                                                                                                                                                       ��������������������������������������������������������������������������    �                                                                                                                                                                                                                       ��������������������������������������������������������������������������    �                                                                                                                                                                                                                       ��������������������������������������������������������������������������    �                                                                                                                                                                                                                       ��������������������������������������������������������������������������    �                                                                                                                                                                                                                       �����                         ��                                    �����    �������������������������� �������������������������������������                                                                                                                                                          ���������������������������������������������������������������������������                                                                              �������������������������� �������������������������������������                                                                                ���������������������������������������������������������������������������                                                                                                                                                                                                                               ���������������������������������������������������������������������������                                                                                                                                                                                                                               ���������������������������������������������������������������������������                                                                                                                                                                                                                               ���������������������������������������������������������������������������                                                                                                                                                                                                                               ���������������������������������������������������������������������������                                                                                                                                                                                                                               ���������������������������������������������������������������������������                                                                                                                                                                                                                               ���������������������������������������������������������������������������                                                                                                                                                                                                                               ���������������������������������������������������������������������������                                                                                                                                                                                                                               ���������������������������������������������������������������������������                                                                                                                                                                                                                               ���������������������������������������������������������������������������                                                                                                                                                                                                                               ���������������������������������������������������������������������������                                                                                                                                                                                                                               ���������������������������������������������������������������������������                                                                                                                                                                                                                               ���������������������������������������������������������������������������                                                                                                                                                                                                                               ���������������������������������������������������������������������������                                                                                                                                                                                                                               ���������������������������������������������������������������������������                                                                                                                                                                                                                               ���                                                                     ��  ����������������������������������������������������������������������                                                                                                                                                        ���������������������������������������������������������������������������                                                                             ����������������������������������������������������������������������                                                                             ���������������������������������������������������������������������������                                                                                                                                                                                                                                 ���������������������������������������������������������������������������                                                                                                                                                                                                                                 ���������������������������������������������������������������������������                                                                                                                                                                                                                                 ���������������������������������������������������������������������������                                                                                                                                                                                                                                 ���������������������������������������������������������������������������                                                                                                                                                                                                                                 ���������������������������������������������������������������������������                                                                                                                                                                                                                                 ���������������������������������������������������������������������������                                                                                                                                                    �                                                                           ���������������������������������������������������������������������������                                                                         ��                                                                                                                                                  ��������������������������������������������������������������������������
�                                                                       P@                                                                       �                                                                           ����������������������������������������������������������������������������                                                                       �@                                                                       H                                                                           ����������������������������������������������������������������������������                                                                       p@                                                                       �                                                                           ���������������������������������������������������������������������������                                                                         ��                                                                                                                                                  ���������������������������������������������������������������������������                                                                                                                                                    �                                                                           ���������������������������������������������������������������������������                                                                                                                                                                                                                                 