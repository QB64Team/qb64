��j  T��                        �    �   0   0 �                                               �    �   0   0 �                                               �    �   0   0 �                                               �    �   0   0 �                                               `  � �0   0 �                                               `  � �0   0 �                                               `  � �0   0 �                                               `  � �0   0 �                                                  � �0   0 �                                                  � �0   0 �                                                  � �0   0 �                                                  � �0   0 �                                               �����;`9ͳ�y��<y�p                                              �����;`9ͳ�y��<y�p                                              �����;`9ͳ�y��<y�p                                              �����;`9ͳ�y��<y�p                                              ��6l ����m��`�0fͳ`                                              ��6l ����m��`�0fͳ`                                              ��6l ����m��`�0fͳ`                                              ��6l ����m��`�0fͳ`                                                                                                                                                                                     o������1���}�0`ͳ`                                                                                                                                                                                                                                                        l������ ͛0`ͳ`                                                                                                                                                                                                                                                       l�6l���`m�6`͛0fͳ`                                                                                                                                                                                                                                                       Ǚ����308�3�}��<y�f�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         �              �                                                   �              �                                                   �              �                                                   �              �                                                  �             �                                                  �             �                                                  �             �                                                  �             �                                                  �             �                                                  �             �                                                  �             �                                                  �             �                                                                                                                                                                                       �             �                                                                                                                    �             �                                                  �             �                                                  �             �                                                  �             �                                                  �             �                                                  �             �                                                  �                                  �              �                                                                              �            ��                   �             �             �            ��                   �             �                                               �              �                                               �              �             �            �                   `             `             �            �                   `             `             �            �                   �             �             �            �                   `             `             @            @                                             @            @                                             �            �                   �             �             @            @                                             >�            >�                   �              �              >�            >�                   �              �              .�            .�                   �             �             .�            .�                                               =�            =�                   �`             �`             �            �                   �`             �`                                              ��             ��                                              �@             �@            ��            ��                   �@            �@            ��            ��                   �@            �@            |�            <�                   l�            l�            <�            <�                   h@            h@             \>             <>                   �            �             ?�             ?�                   ��            ��             �2             �2                    l�             l�             L2             ,2                    l�             l�             D>             t>                   �            �             ��             W�                   ��            ��             �             �                   �             �              T             D                   �             �             �4            �4                   �            �            k�            ��                   ��             ��            �            �                   a             a             �            �                   a              a             J�             �                   !�            �             ��             ��                   ��            ��            Ύ            Ύ                    �            `�            �             ��                   ��             �            
3            γ                   )�            �            ��            O�                   ��            ��            �-            �-                   h@            H@            I�            !                   �                          �            �                   �            ŀ            �            �                   �            G�            �                               D�            ��                                           ��            �            (            �                   A             �             ^            �                   �             �             :            8                   �                          d                                                         (             :                    0�             �             ^             >                    /�             
�             x             p                    9�                           &             0                                                jP             ~�                                                v�             ~�                    o�                           ^�             H`                    1              :              HH             H`                    ^�                           �             T                    !              ~              x             
\                    _              z              <�             <�                    c              4              �             @                    <              0              �             �                    �              .              -x             �                    �              *              9�             9�                    �              t              �             �                    X                            �@            ��                    @              \             ��            ��                   �              T             {�            !�                    �              �             !             !�                   z              @              R�             9P                    �             �              5�             )p                   |             �              �             �                   �              �              F@             !                     �              �              B�             s�                                 �              ��             S�                   �              �              �             �                    �             �              R`             C                    `              �             �             �@                                 p             k�            ��                   �             P             �@            �                                 �             ��            �                    �                           J              �@                                �              ׀             ��                   �             �             ΀            �                    0             @                           �                    �                           
             ΀                                 �             ׀            O�                   �             �             �             �                    `             @             I�                                �                           �             �                                  �             �             �                    �             @             �                                 @             �                                              �                           (                                 (@             ?�             	�             	�                    7�             >�             :             8                    �                           	d             	                                                h             z                    0�             ;�             �             �                    ?�             :�             x             p                    9�             =              f             p                    6              8              0             4                                                �             �                    �                           $                                  i              j              (                                  
�                           8             <                    �              �              *�             
�                                                                                 {              z              2             
                                                >             >                    ��             ��             -�             �                    ��             ��             9             9                    q              1                                               q              1              )             {                    Y�             Y�             Z�             {�                   ��             W�             {O             !O                    �@             �@             !O             !O                   P@             @             R��            9�                   ��            ��             ���            )�                  �            ��             s��            s��                  �p             �p             �o�            !/�                   �`             �`             B�@            s�@                  �             ��             ���            S��                  ��             ��             �@            �@                  �p            �p             Ro@            C@                  b`             �`             ��           �D�                  �            q�            kĀ           �Ā                  ��            Q�            �G�            ��                  `            �`             ���            ��                  �`            `            J             �A                   �            ��            ׁ             ��                   ��            ��            ΃            �                   0@            @@                         �                   �@             @            
             ΀                                 �             ׀            O�                   �             �             �             �                    `             @             I�                                �                           �             �                                  �             �             �                    �             @             �                                 @             �                                              �                           (             �                    @             �             ^             �                    �             �             :             8                    �                           d                                                             (             :                    0�             �             ^             >                    /�             
�             x             p                    9�                           &             0                                                
P             �                                                �             �                    o�                           �             `                    1              :              H             `                    ^�                           �             T                    !              ~              -x             
\                    _              z              �             �                    c              4              1�             @                    <              0              �             �                    �              .              -x             �                    �              *              9�             9�                    �              t              �             �                    X                             )@             {�                    @              \              Z�             {�                   �              T              {�             !�                    �              �              !              !�                   z              @              R�             9P                    �             �              ��             )p                   |             �              s�             s�                   �              �              �@             !                     �              �              B�             s�                                 �              ��             S�                   �              �              �             �                    �             �              R`             C                    `              �              �             �@                                 p             k�            ��                   �             P             �@             �                                 �              ��             �                    �                           J              �@                                �             ׀             ��                   �             �             ΀            �                    0             @                           �                    �                           
             ΀                                 �             ׀            O�                   �             �             �             �                    `             @             I�                                �                           �             �                                  �             �             �                    �             @             �                                 @             �                                              �                           (             �                    @             �             ^             �                    �             �             :             8                    �                           d                                                             (             :                    0�             �             ^             >                    /�             
�             x             p                    9�                           &             0                                                
P             �                                                �             �                    o�                           �             `                    1              :              H             `                    ^�                           �             T                    !              ~              -x             
\                    _              z              �             �                    c              4              1�             @                    <              0              �             �                    �              .              -x             �                    �              *              9�             9�                    �              t              �             �                    X                             )@             {�                   @             \              Z�             {�                   �             T              {�             !�                    �              �              !              !�                    z              @              R�             9P                                x              ��             )p                   �             �              s�             s�                                  P              �@             !                     p              @              B�             s�                   �             �              ��             S�                   �             �              �             �                                                 R`             C                                                   �             �@                   `             p             k�            ��                   3�             3�             �@             �                                                ��             �                                                J              �@                                             ׀             ��                   9�             9�             ΀            �                                                              �                                                  
             ΀                                             ׀            O�                   <�             <�             �             �                                                I�                                                              �             �                    q�             Q�             �             �                    �p             �p             �                                                                                                                            (             �                    8�             8�             ^             �                    �0             �0             :             8                    �             �             d                                                               (             :                    0             0             ^             >                    ��             ��             x             p                                                &             0                                                  
P             �                   �             F              �             �                   9�            9�             �             `                    @              @              H             `                    �                             �             T                    �              �              -x             
\                   ��            ��             �             �                    b              b              1�             @                                                  �             �                    p�             p�             -x             �                   ��            ��             9�             9�                                                �             �                                                  )@             {�                                              Z�             {�                   �             �              {�             !�                                                !              !�                                                 R�             9P                   �             �              ��             )p                   s             s              s�             s�                   �             �              �@             !                                                   B�             s�                   �             �              ��             S�                   ?             ?              �             �                     @              @              R`             C                                                   �             �@                   `             `             k�            ��                   3�             3�             �@             �                                                 ��             �                                                 J              �@                   0             0             ׀             ��                   9�             9�             ΀            �                                                              �                                                  
             ΀                                             ׀            O�                   <�             <�             �             �                                                I�                                                              �             �                    �             �             �             �                    >p             >p             �                                                                                                                              (             �                     �              �             ^             �                    ?0             ?0             :             8                     �              �             d                                                               (             :                    `0              0             ^             >                    _�             /�             x             p                    p                            &             0                                                  
P             �                                   X              �             �                    ��             _�             �             `                    `              8              H             `                    �                            �             T                    @              4              -x             
\                    ��             ��             �             �                    �              |              1�             @                    |              0              �             �                   �              �              -x             �                                 �              9�             9�                   �              t              �             �                    �              0              )@             {�                    �             x              Z�             {�                                p              {�             !�                   �              �              !              !�                   �              `              R�             9P                                 �              ��             )p                   �             �              s�             s�                                �              �@             !                    �              �              B�             s�                                �              ��             S�                   �             �              �             �                                 �              R`             C                    �              �              �             �@                                 �             k�            ��                   �             �             �@             �                                 �              ��             �                    �             �             J              �@                                @             ׀             ��                   �                           ΀            �                    8             �                           �                    �                           
             ΀                                �             ׀            O�                   �             �             �             �                    p             @             I�                                �                           �             �                                  �             �             �                    7�                           �                                 `             �                                              /�                           (             �                                                ^             �                    /�             ,              :             8                    0�             �             d                                                             (             :                    `@             /�             ^             >                    _�             .�             x             p                    q�                           &             0                    .                            
P             �                                   ^              �             �                    ��             \              �             `                    a�             ;              H             `                    �@                           �             T                    @�             4              -x             
\                    ��             �              �             �                    À             ~              1�             @                    |              0              �             �                   �              �              -x             �                                 �              9�             9�                   �              t              �             �                    �              0              )@             {�                    �             x              Z�             {�                                p              {�             !�                   �              �              !              !�                   �              `              R�             9P                                 �              ��             )p                   �             �              s�             s�                                �              �@             !                    �              �              B�             s�                                �              ��             S�                   �             �              �             �                                 �              R`             C                    �              �              �             �@                                 �             k�            ��                   �             �             �@             �                                 �              ��             �                    �             �             J              �@                                @             ׀             ��                   �                           ΀            �                    8             �                           �                    �                           
             ΀                                �             ׀            O�                   �             �             �             �                    p             @             I�                                �                           �             �                                  �             �             �                    7�                           �                                 `             �                                              /�                           (             �                                                ^             �                    /�             ,              :             8                    0�             �             d                                                             <(             ?:                    `@             /�             ;^             =>                    _�             .�             x             p                    q�                           &             0                    .                            ~P             ~�                                   ^              ~�             ~�                    ��             \              �              `                    a�             ;               H              `                    �@                           ��             �T                    @�             4              �x             �\                    ��             �              8�             8�                    À             ~              9�             8@                    |              0             8��            8��                   �              �             ;��            ;��                                 �              8              8                    �              t              8             8                     �              0             D�             D�0                   �             �             ��            ��                   �             �              8              8                                                8              8                                                �}�            �}�                   �             �             ���            ���                   �             �             8�            8�                   �              �             8�            8�                    �              �             �=�            �=�                   �             �             ���            ���                   �             �             8�            8�                   �              �             8�            8�                   �              �             ��            ��                   �             �             ���            ���                   �             �             8�            8�                   �             �             8�            8�                   
�              �             D             D                    �             �             ��            ��                   �             �                                                                                                                                              8�            8�                                �             ;��            ;��                   �             �                                                  0             �                                                  �             �                                                                 �                                                  �             @                                                  `             �                                                  �                                                                                                                                  �                                                                 �             �                                                                                                                    @             �                                                  �             �                                                  �                                                                                                                                                 �                                                  �                                                                                                                                   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               <    �0      <    �             �`     �0   �`     �                                                                                                                                                                                                              f     �      f     �              `      �    `      �                                                                                                                                                                                                              `     �      `                   `      �    `                                                                                                                                                                                                                    `�����7�     `����9���         g�<y�||�7�  g�<y�||9���                                                                                                                                                                                                          <͛�l���l     <͛�l��6�0         3l�f͛v���l  3l�f͛v��6�0                                                                                                                                                                                                          ͛6o��l     ͛6o��6��         ?o�`͛f��l  ?o�`͛f��6��                                                                                                                                                                                                          ͛6l�l     ͛6l�6�          0l`͛f��l  0l`͛f��6�                                                                                                                                                                                                           f͛6l��l     f͛6l�ٳ6�0         3l�f͛f��l  3l�f͛f�ٳ6�0                                                                                                                                                                                                          <��3��f     <��3������         g�<y�f|�f  g�<y�f|�����                                                                                                                                                                                                           �  `           �  `                     �            �                                                                                                                                                                                                                  � �           � �                     � �           � �                                                                         