��d   ��?                          �                                                                                                   �                                                                                                  �                                                                                                  �                                                                                                  �                                               @                                                �                                               @                                                �                                               �                                                �                                               �                                             >  �                                              F                                             >  �                                              F                                               �                                                                                             �                                                                                           �� �                                                                                           �� �                                                                                          ��  �                                              
1                                            ��  �                                              
1                                            ��p                                               "                                            ��p                                               "                                            ��   �                                           $                                           ��   �                                          <$                                           ���׀�                                            (h                                           ���׀�                                           ���h                                           ���� ?�                                            (���                                          ���� ?�                                            ?�����                                           ���+ �                                           ^4��                                            ��� �                                           ���                                            � p �                                          �?t��                                            �   }�                                          ����                                            >    �                          ��������������  �?8$��                          ��������������   >    |�                                          �?8��                          �������������   �  �                          �              '�>8D��                         �               �  |�                          �������������  '�>8D��                         �������������   � �                          �              7�L?���                         �               �  �                          �������������  7�L8���                         �������������    � ��                          �              ����                           �                `  ?�                          �������������  ��p@                           p            p    � ��                          �������������� �Q����                           ��������������    � �                          p            p �ќ��                            p            p    � ��                          �������������� ���8���                           ��������������    � ��                          p            p ���8���`                          p            p  �    p                          ��������������  ����?�                          ��������������  �     p                          p            p  ����9�                          p            p �     �                          ��������������  ��87                           �������������� �      �                          p            p  �`�87�                          p            p � ?�   <                          ��������������  ��0�                           �������������� �     <                          p            p  O�Dy0�<                          p            p ��?�                            ��������������  ����                           �            � � 
                             p���   ����p J��                          p            p ��?�  �                          ��������������  �����                           �            � �    �                          r6�m�$�I#m��rp �}��                          p            p ��   �                          ��������������  �����%?                          �            � �@    �                          p���   ����p �O����%?                          p            p  �   �                          �������������� �w��� �                         �            �        �                          p���   ����p ����"�                         p            p  �    À                         ��������������  ?����e0                          �            �       À                         r6�m�$�I#m��rp ?���e3�                         p            p     8 ��                         ��������������  ?�����p|                          �            �       ��                         p���   ����p ?�����p}�                         p            p     | �                         ��������������  �����x�                          �            �       �                         p���   ����p �����x��                         p            p 8   8|   �                         �������������� �������                          �            � 8   8   �                         r6�m�$�I#m��rp ;��������                         p            p 8   ||  �                         �������������� ������                          �            � 8   |   �                         p���   ����p ;�������                         p     �     p p ��8  8p                         ������������� ��}> �                          �     �     � p ��   8p                         p��� �����p q��} �p                         p     @     p p �� �p                         ������ϟ������  ?��)���                           �     ?�     � p   �   p                         r6�m�$��#m��rp p>�)��< p                         p     ;�     p p �� � p                         �������O������  ������                          �     �     � p  �    p                         p��� �����p p����p                         p     k�     p � �| � x                         �������/������  �������                          �     w�     � �  |  � x                         p��� �����p �������x                         p     P(     p   �8 � 8                         �������������?�������                          �     ��     �   �8 � 8                         r6�m�$��#m��rp�?�������8                         p     �     p � �  � 8                         ������/����������������                         �     �x     � � 	    � 8                         p��� ������p���������                         p     ��     p � �  �                          ������?������� ���������                         �     �     � �                                 p��� ������p���<�����                         p     �(     p � � �                          ������?������� ��|����                           �     �     � � �                              r6�m�$�y#m��rp���|���> 8                         p     �8     p�    :>                           ������?������� ������{�$                         �     �8     � �    >                           p��� �8����p�������{�<                         p      p     p�     <                         �������������� ��x�o�                         �     `0     � �     8                         p��� `p����p���h�o�<                         p     �     p�8   �� <                         �������������� ��� N    ��������             �     pp     � �8   �� 8    ��������             r6�m�$��#m��rp���� N<                         p     �     p�� �� <    ��������             ������������� o����           �            �     ?�     � �   �� 8           �            p��� ?�����p�o�<���    ��������             p           p� � �� >   ���������            ������������� �����"  �           @            �     �     � �    �� 8           @            p��� �����p�����"  �   ���������            p            p� � �� ~   ���������            ������������������                          �            � �    �� x                        r6�m�$�I#m��rp��O�� ~   ���������            p            p� �p�� v   �      �            ���������������O����A�   �������            �            � p  � �� x   �������            p���   ����p�O����]�~   �      �            p            p������ v          �            ���������������~���  �   ��������            �            � p�  �� x   ��������            p���   ����p�yO� �~          �            p            p������ v   �       �            ���������������8��,"�   !�������            �            � p�  �� x   !�������            r6�m�$�I#m��rp�8'$"�~   �       �            p            p������ �   =�       |            ���������������9��> @   B��������            �            � 8� P�� �   B��������            p���   ����p�9<u" @�   =�       |            p            p�� p�� �   {�       >            ���������������`?�|, p    ���������            �            � 8�   �� �   ���������            p���   ����p�`?�,$ p �   {�       >            p            p��    �   �                    ���������������D?� �x   ����������           �            � �    �  �      ��           u�$�H�m�ܒI$�p�D?� �x!�   �[m�$�H�l            p            p�     > �  �        �           ���������������;�� ��  ���������@           �            �      > �         �@           w�  ����   p�?�� ���  ����  ���           p            p�       �  �        �           ���������������;��#��   #���������            �            �        �  "        �            w�  ����   p�;��#���  ����  ���           p            p�       �  �        �           ���������������#��#�    G���������           �            �        �  D        |           u�$�H�m�ܒI$�p�#��#� �  ��m�$�H�m��           p            p��       p        �           ����������������� �   ����������           �            � �      �  �        >           w�  ����   p���� o��  w���  ����           p            p��        �         �           ����������������(�   !���������           �            � �      �  !                   w�  ����   p���(��  ����  ����           p            p�� �     =�         |           ���������������)��   B?����������           �            � � �   �  B         �           u�$�H�m�ܒI$�p��)���  =��m�$�H�m�|           p            p�� �   <  {�         >           ���������������  	#�   �����������           �            � � �   ?�  �@        �           w�  ����   p�� 	+�?�  {����  ���>           p            p�� �   �  �                     ���������������� 	7�  ������������          �            �  x �   �� �        ��          w�  ����   p�� 	7���  ����  ���           p            p�� �  � �          �          ���������������� 	7   �����������@          �            �  | �  ��          �@          u�$�H�m�ܒI$�p�� 	7�� ��m�$�H�m��          p            p �� �  �8 �          �          �������������� ��    8 #�����������           �            �  > �  �� "          �           w�  ����   p ��  �� �����  ����          p            p �� �  �8 �          �          �������������� ��    8 G�����������          �            �   �  �� D          |          w�  ����   p ��  �� �����  �����          p            p ����   8 p          �          �������������� ��    8 ������������          �            �  ��  �� �          >          u�$�H�m�ܒI$�p ��� �� u��m�$�H�m���          p            p ��    | p �           �          �������������� �    p !�����������          �            �  �    �� !                    w�  ����   p �� �� �����  �����          �            x ��    � � =�           |         ������������� �     � B?������������                     �  �    ��  B           �          ��  ����   x ��  ��� =�����  ����|         �            | �~   � � {�           >         ������������� �      � �������������                     �  �   ��  �@          �         ��$�H�m�ܒI$�| ��  ��� {���m�$�H�m��>         �            > ?��   � �                     ������������� ?�      ���������������                    �  ��  �� �          ��        �  ����   > ?���  ��� �����  ����         �             ?��  ��            �        ?��������������?�     ��������������@        8            ��  ��  ��            �@        ǀ  ����    ?���  ��������  �����        �            �?�����<��            �        �������������@?��    <�#�������������         x            �@  ����� "            �         ��$�H�m�ܒI$��?��������܍��m�$�H�m���                     ���������            �         �������������� ��    ��G�������������         �            �  ����� D            |        �  ����   ���������������  �����        >             �������p            �        A���������������   ����������������        A�            |  �����?� �            >        >�  ����   �����������p����  �����        |             ����   ��             �        ������������������   �!�������������        ��            >  x����� !                    |�$�H�m�ܒI$������������䍶�m�$�H�m�܀�        �              ���� �  =�             |       ����������������� �  B?��������������       �              > ���� B             �        �?�  ����   ���������� =�����  ���� |       �              |����� ? {�             >       �������������������� ? ���������������       �            �  �  �� �@            �       ��  ����   �|�������� {�����  ���� >       �              >�� ��  ~ �                     ����������������� ��  ~����������������                   �  � ����            ��      �m�$�H�m�ܒI$��>�������� �$���m�$�H�m�ܐ       �              ��     ��              �      ?������������������     ����������������@      >             �� �����              �@      ���  ����   ���������� ����  ���� �      �              ���    ��              �      ���������������@��    �#���������������       |             �@ ����� "              �       ���  ����   ����������� ����  ���� �                     ���    ��              �       ���������������� ��    �G���������������       �              �   ����� D              |      m�$�H�m�ܒI$������������$���m�$�H�m�ܒ�      >               ���   �p              �      A������������������   �����������������      A�              |  ?���� �              >      >��  ����   ����������p ����  ���� �      |               �?��   ?��               �      �����������������?��   ?�!���������������      ��              >  ���� !                    |��  ����   ���?�������� ����  ����  �      �                ���  ��=�               |     ������������������  ��B?����������������     �                ���  B               �      �$�6�m�$�I#m��rI ��������=��rI$�6�m�$�I#m�|     �                |��� � {�               >     �������������������� � �����������������     �              �   ��  �@              �     �  ���   ����  |������ {���   ���   ��>     �                >��� �� �                     �������������������� ��������������������                   �   �  �              ��    �  ���   ����  >������ ���   ���   ��     �                �������                �    ?�����������������������������������������@    >               ��                     �@    �$�6�m�$�I#m��rI$��������rI$�6�m�$�I#m��    �                �������                �    �����������������@�����#�����������������     |               �@      "                �     �  ���   ����  ����������   ���   ���                     �?������                �     ������������������ ?�����G�����������������     �     ?�����     �       D     �����     |       ���    ���  �?���������          ����    >      ?�����     ������p     �����     �    A�������    ������������������    ������    A�     @         |      �               >    >	$�6�m�������rI$�������u��rI$�������I#m���    |      �����     ����� �     ?�����      �    ��������    ���������� !������    ������    ��     �         >      !     @             |   ����������  ����� ����  ?�����  ����    �      ������      � ��� =�     �����      |   ������     ������ ��� B?������    �������   �                    B      �         �    �   �����������   � ��� =����  �����  ���|   �     �    |      | ��� {�     �    >      >   ������������������ ��� ������������������   �    �����     �      �@    �����     �   �I$�6�m�    }��rI$�| ��� {���rI$�    >�I#m��>   �     �    >      >  ��  �     �             ������������������  �� �������������������       �����     �     �    ������    ��  �   ���    >���   >  ��  ���� �      ���   �     �               �     �    �     �  ?������/�����������������������������������@  >     /������    �������     �����@    �@  �   ���    ��        ����� �    � ����  �     �    �     �������     �    �     �  ������O�����������      #������'�����?������   |     O�����@    �      "     '�����      �   �I$�6�o�    ��rI$��������m��rI'�    �I#m���        p    �     �������     �    �     �   �������������?������      G������G�����������   �      ������      �      D     G�����     |      ��p    ���   ����������� �    � �����  >      >�    �     ������p     x    �     �  A������������������      �������������������  A�     A�����     |      �      ������     >  >    ���    ���   ������w���� x    � �����  |      }�    �            �     >�     �      �  ������������������������������������������  ��     ������     ?������     A�����       |I$�6�}�    ��rI$�       �m��rI>�     �I#m��`�  �      ��     �            �     }�     |      | �����������������������?������������������� �    �����     ������      �������     �  �    ���     ���   `      ����� }�     | ����| �     ��     |            �     ��     >      > ������������������������������������������ �    ������     ������@    ������     � �`   ���     }��   p      ����� ��     > ����> �     ��     >                 ��            ��������������������������������������������     ������     �������    �������    ���rI$�6���     >�rI$�0      #m��rI��     I#m��p �     ��   �                  ��   p �     �?������ �����������������������������������@>      �������    ������     ������@    �@��   ���     �   |      ������     �������     ��  � �                ��   � �     �������@���������������������� �����?������ |     @������@                 ������      � ��   ��     ��   ���   ������     ������      �  � �                ��  � �     � �����������G��?�����������������@���#�������� �      �������                 @������     |rI$�6��  @ �rI$�6�m�$�I#m��rO��    �#m��r�>      >��  � �                �  � �     �A������� ���������������������������S��������A�     A ������                 �������     >>�   ���  � ��   ���   �����  q ������|      }��  � �                >��  �  �      ��������� ���G�������������������  ���#����������     � ?������                A ������     |�   }��F ��   ���   ����>��#  ����� �x      ���  �  �                }��� �  |      x�������  ����������������������  ��������������     ������                � ?�������     �xrI$�6���  �rI$�6�m�$�I#m��r}��  }#m��r@xp     ���� �  |                ����  �  >      8�������  ���������������������  ?�����������ď�     ��������                �������     �p�   }��   }�   ���   �������  >���� 8p     ����  �  >               ���� p        8�������  ?���������������������  ������������ď     ��������                ����x����    �p��   {�� 
1  >�   ���   ������ �  ���� 8p     ����p                   ����8    �     8�������  ?���������������������� �����������Ď      ���������               ��������@    �p�rI$�7��"  rI$�6�m�$�I#m��s��
  �m��rH8p     ����   ��              ����  ��     8�������@ ?�������������������� ����?�?�����Č     @��������@                ��������      �s��   o��<$ �   ���   ������ ����� 8p     ����׀��              ���������     8��������  >(�?�?���������������@  ?�������Ĉ      ��������               @��������     Dw��   _����h �   ���   ��������4 ����� 8p     >������ ?��              �������     8�������   (��������������������  �O������Ĉ     A ���� ?��               � ������     Dq$���m��� ?�������m�$�H�m�ܒI$�� ����@��I$���p     }�����+ ��              >�����?� �     8�������  ^4������������������  �/�������Ĉ     �  ��� ��              A  ���?��     Dp ���}�� ��� �����  ����   >���?���  �   ��p     ���� p � �              }��?� 8 ?� |     8������ �?t������������������ ��:ć�������Ĉ      �   }��              �  ?�   >���     Dp ����������  �����  ����   }����ŀ |   ��p    ���>    � |              ���   ?� >     8������ �?8$������������������ ��?�G�������Ĉ      >    |���                   >��     Dq$���m����?8�� }��m�$�H�m�ܒI$�����?�� >�I$���p    ����  � >             ��� �  ?�      8������ '�>8D����������������� �"?��������Ĉ      �  |��                �  >x?��    Dp �������>8D��>����  ����  ����"?���   ��p    ���� �              ���� �� �    8������  7�L?������������������ �&�G������Ĉ       �  ���              �  ?���@    Dp �������L8������  ����  ����&D@@�  ��p    ��� � �� �            ��� � �� �    8������@ �������������������  �L�?���?����Ĉ    @   `  ?���@                �  ���     Dq$���o�����p@  ��m�$�H�m�ܒI'�����8   �I$���p    �  � �� �            ��  � �� �    8��������Q����?��?�������������@���T�������Ĉ     �   � ���             @   �  ����    Dp �����ќ��   ����  ����  �����Tx�  �  ��p    >��  � �� �            �   � �� �    8������ ���8���������������������oH��������Ĉ    A    � ����             �    � ����    Dp ��������8���` ����  ����  ���oL��0 �  ��p    }���    p �            >���   �8  �    8������  ����?����������������  ��Ο��������Ĉ    �  �     ��            A  p     �?��    Dq$���}������9� ��m�$�H�m�ܒI>����x�Μ��  �I$���p    ����     �  �            }��� �   x  |    8�����  ��87���������������  �?����������Ĉ    �      ���            �  �      ���    Dp ������`�87�  ����  ����  }���0|��  |  ��p   ���� ?�   <  |            ���� �     >    8�����  ��0����������������  �?��g�������Ĉ    �     ?���             �     ���    Dp �����O�Dy0�<  }���  ����  ���'�"<�g  >  ��p   �����?�    >           ����p�  �      8�����  �������������������  ����� �������Ĉ    � 
   ���            �    �����   Dq$������J��  >�m�$�H�m�ܒI�����?��  I$���p   �����?�  �             ������  �  �   8�����   ��������������������  ����?� ������Ĉ     �    �����           �    ����@   Dp ������}��  ��  ���� �����>�?�  � ��p   �����   �  �          ������  �  �   8�����@  �����%?��������������   ���������?���Ĉ   @ �@    ����@            �     ���    Dp �����O����%?  ���  ���� ����'����� � ��p   ���   �  �          ��� �   �  �   8������ �w��� ���?�����������@ ���� ������Ĉ    �        ���?�����������@        �?��   Dq$���������"� �          ����C���� �$���p   ��� �    À �������������� p    �� �   8�����  ?����e0��            � ����2�?�����Ĉ   !        ����            �       ����   Dp �����?���e3� ������������������2�� � ��p   ���    8 �� ���������������     ��  �   8�����   ?�����p|?��             �����8>�����Ĉ   "  <      ����                   ����   Dp �����?�����p}� ��������������������8>�  � ��p   ���    | �  ���������������    > ��  �   8�����  @�����x���              �����<�����Ĉ   "  \      ���             .      ����   Dq$�����������x��  ��������������������<�  �$���p   ��8   8|   �             ���   >   p  �   8�����  ����������������������  A�����ÿ�������Ĉ   "  �   8   ���������������  \      ��   Dp ����;��������             ��������˿��  � ��p   ��8   ||  �             ��   >>  p  �   8����� ��������������������  �����?��������Ĉ   " 8   |   ���������������  �   >   w��   Dp ����;�������             ���������p  � ��p   ��p ��8  8p             ��8 �  8  �   8����� ��}> ���������������  �澈 �����Ĉ   " p ��   8s�������������� 8 @   ;��   Dq$�����q��} �p             ��8�f>� 8  �$���p   ��p �� �p             ��8 �  �8  �   8�����  ?��)��� ��������������  ����� �����Ĉ   " p   �   q�������������� 8      9��   Dp ����p>�)��< p             ��8d��� 8  � ��p   ��p �� � p             ��8 � � 8  �   8�����  ������ ��������������  ������ �����Ĉ   " p  �    p�������������� 8     8��   Dp ����p����p             ��8�����8  � ��p   ��� �| � x             ��x�> � <  �   8�����  ������� �������������  ������� ����Ĉ   " �  |  � x������������� x �>  @ <�   Dq$������������x             ��x�����G�<  �$���p   ��  �8 � 8             ��  � �   �   8����� !�?������� ?������������� ���~���� ?����Ĉ   "    �8 � 8?�������������   @  � ?�   Dp �����?�������8             ����������  � ��p   ��� �  � 8             ��p �  �   �   8����� C���������������������� !��������������Ĉ   " @� 	    � 8�������������  p �   @ �   Dp �������������             ���������G��  � ��p   � � �  �              ��p �  �   �   8����� � ���������������������� A ��g���������Ĉ   " ��        ������������� @p        �   Dq$�������<�����             ��p�g����  �$���p   � � � �              � p �  �   �   8����� ��|����  ������������� � {d�G��� ����Ĉ   " � �     ������������� �p @     �   Dp ������|���> 8             �p{�>G��   � ��p   ��    :>               � �        �   8����� ������{�$������������� �C��D��=�����Ĉ   " �    >  ������������� p      �   Dp ����������{�<             � �C��D��=�  � ��p   ��     <             � �   ��   �   8����� ��x�o�������������� ���<@7�����Ĉ   " �     8������������� p   �� �   Dv�rI����h�o�<             � ���4@7�  ��rI8p   ��8   �� <             � �   �   �   8����� ��� N ������������� ���΀'� ����Ĉ   " �8   �� 8 ������������� p   �  �   Dw�� ����� N<             � ���΀'�  ��� 8p   ��� �� <             � � �  ��   �   8����� o���� ������������ �7��� � ���Ĉ   " �   �� 8 ������������ p    ��     Dw�� ��o�<���             � �7��@�  ��� 8p   �� � �� >             �� � ��   �   8�����  �����"  � ?�������������w���~  C ?���Ĉ   "  �    �� 8 ?������������ p    ��  ?   Dv�rI������"  �             ��w��~  _  ��rI8p   �� � �� ~             �� � �� ?  �   8�����@����   ������������ ���_�~   ���Ĉ   "@ �    �� x ������������  x    �� <    Dw�� ���O�� ~             ������� ?  ��� 8p    � �p�� v             �� �8�� ;  �   8������O����A� ������������@�'���� �� ���Ĉ   "� p  � �� x ������������@ 8  @ �� <    Dw��  �O����]�~             ��'�G��.��?  ��� 8p    ������ v              ���|�� ;  �   8����� �~���  � ��������������?_��  ` ���Ĉ   #  p�  �� x ������������� 8�  �� <    Dv�rI �yO� �~              �<��� `?  ��rI8p    ������ v              ���|�� ;  �   8����� �8��,"� ������������ ����� ���Ĉ   "  p�  �� x ������������  8� �� <    Dw��  �8'$"�~              ����?  ��� 8p    ������ �               ���|�� s  �   8����� �9��> @ ������������ ���n�  ���Ĉ   "  8� P�� � ������������  � ( �� |    Dw��  �9<u" @�               ��:�   ��� 8p    �� p�� �               �� 8� s  �   8����� �`?�|, p   ������������ �0�> 8 ���Ĉ   "  8�   �� �  ������������  �  � |    Dv�rI �`?�,$ p �               �0� 8  ��rI8p    ��    �               ��   ?� �  �   8����� �D?� �x                �"��@< ���Ĉ   "  �    �                �   ?� �    Dw��  �D?� �x!�               �"��@<�  ��� 8p    �     > �               �       �  �   8����� �;�� ��               ���`� ���Ĉ   "       > �                       �    Dw��  �?�� ���               ���`��  ��� 8p    �       �               �       �  �   8����� �;��#��                �����  ���Ĉ   "         �                       �    Dv�rI �;��#���               ������  ��rI8p    �       �               �       �  �   8����� �#��#�                 �����  ���Ĉ   "         �                       �    Dw��  �#��#� �               ������  ��� 8p    ��                    ��     �  �   8����� ��� �                ���?�  ���Ĉ   "  �      �                �      �    Dw��  ���� o��               ����7��  ��� 8p    ��                     ��        �   8����� ��(�                �~?�  ���Ĉ   "  �      �                �      �    Dv�rI ���(��               ��~?��  ��rI8p    �� �                   �� �     �   8����� �)��                 ���  ���Ĉ   "  � �   �                � �   �    Dw��  ��)���                �����  ��� 8p    �� �   <                �� �     �   8����� �  	#�                 �  ��  ���Ĉ   "  � �   ?�                 � �   �    Dw��  �� 	+�?�                �� ���  ��� 8p    �� �   �                �� �   x  �   8����� �� 	7�                 �� ��  ���Ĉ   "   x �   ��                 < �   �    Dv�rI �� 	7���                �� ���  ��rI8p    �� �  �                �� �   �  �   8����� �� 	7                  �� ���   ���Ĉ   "   | �  ��                 > �   ��    Dw��  �� 	7��                �� ��� ��  ��� 8p     �� �  �8                � �  �  �   8�����  ��    8                �     ���Ĉ   "   > �  ��                  �  ��    Dw��   ��  ��                �  ��  ��� 8p     �� �  �8                ���  �  �   8�����  ��    8  ������������  �  
   ���Ĉ   "    �  ��  ������������   ��  ��    Dv�rI  ��  ��                �� 
��  ��rI8p     ����   8  ������������  ���  �  �   8�����  ��    8              �  �   ���Ĉ   "   ��  ��               ��  ��    Dw��   ��� ��  ������������  �� ���  ��� 8p     ��    | p ������������  ?��    > 8  �   8�����  �    p              ?�  	  8 ���Ĉ   "   �    ��               �    ?��    Dw��   �� �� ������������  ?�� 	?��  ��� 8p     ��    � � ������������  ?�|    | x �   8�����  �     �             � ?�     x ���Ĉ   !   �    ��              �  �    ��    Dv�rI  ��  ��� ������������  ?��  �� ��rI8p     �~   � � �          � ?�?   � x �   8������ �      � ?�����������@ ?�      x ���Ĉ    �  �   ��  ?�����������@  �   ���    Dw��   ��  ��� �          � ?��  ��� ��� 8p   � ?��   � �          � ��  ?� � �   8�����@ ?�      � �����������  �       � ?���Ĉ   0@  ��  ��  �����������   ��  ?��  0   Dw�� � ?���  ��� �          � ���  ?��� ��� 8p   � ?��  � @          � ���  ?��� �   8�����  ?�     �  ������������ ��    �� _���Ĉ   8    ��  ��   ������������   �  ?�  P   Dv�rI� ?���  ��� @          � ���  ?��� ��rI8p   � ?�����<� >�          � ������ `   8����� ?��    <� A?����������� ��    �  ����Ĉ   <   �����  A?�����������   �����   �   Dw�� � ?�������� >�          � �������� o�� 8p   � ������� }�           � �|?���|� >�   8����� ��    �� �?����������� �|    |� A���Ĉ   >  �����  �?�����������   �������  A   Dw�� � ��������� }�           � ��������� >��� 8p    � ������ ��           | ������� }�   8����� �   �������������� ��   �� �?���Ĉ      �����?� @          �   p�����  �    Dq$���� ��������� ��m�$�H�m�ܒ@| ��������� }�$���p    | ���   ��            > ���  ?�� ��   8������ ���   �������������� ���  ?�����Ĉ   �   x����� �          �   <���� @   Dp ��| ������������  ����  > ��������� �� ��p    > ��� �  �             ����� ��    8������ ��� �  ������������������� �����Ĉ   �   > ����            ��   ��� �   Dp ��> �������� ����  ����   ����������  ��p     ����� ? �            ������ ��    8������������ ? #�������������@����� �����Ĉ   ��  �  �� "           �@  �  ?��     Dq$��� �������� ��m�$�H�m�ܒH�����������I$���p    ��� ��  ~ �            ��� �  ? �    8������@�� ��  ~ G������������� �� �  ? #����Ĉ   �@  � ��� D            �   ����� "    Dp ����������� ����  ����  ��������� �  ��p    ���     � p            � ��     ~ �    8������ ��     �  �������������� ��     ~ G����Ĉ    �   �����   �            |  ������ D    Dp ����������� w���  ����  � �������� �  ��p    � ��    � >�            � �    � p    8������ ��    � A������������� �    �  �����Ĉ    |  �����  A            >   �����   �    Dq$���� �������� >��m�$�H�m�ܒI� ������� rI$���p    � ��    � }�             � ��   � >�    8������ ��    � �?������������� ��   � A����Ĉ    >   �����  �                ����  A    Dp ���� �������� }����  ����   � ������� >�  ��p     � ��   � ��             | ?��   � }�    8������ ��   ��������������� ?��   � �?����Ĉ       ?���� @            �   ����  �     Dp ���� ������� �����  ����   | ?������� }�  ��p     | ?��   ?��              > ��   � ��    8������� ?��   ?���������������� ��   �����Ĉ    �   ���� �            �   ���� @    Dq$���`| ?��������6�m�$�H�m�ܒI > ������� ��I$���p     > ��  ���               ��   ���     8������� ��  ��������������������   �������Ĉ    �   ���               ��  ���  �    Dp ���> ������������  ����    ��������   ��p      ��� � �              ���� ���     8����������� � #���������������@��� �������Ĉ    ��   ��  "             �@   ?��       Dp ��� ������ �����  ����   ���������   ��p     ���� �� �              ���� � �     8�������@��� �� G��������������� ��� � #�����Ĉ    �@   �   D              �    ��  "     Dq$���l������� ���m�$�H�m�ܒI$������� ܒI$���p     ������� p              � ������ �     8������� ������  ���������������� ������ G�����Ĉ     �          �              |        D     Dp ���������� w����  ����   � ������ �   ��p     � ����� >�              � ?����� p     8������� ����� A��������������� ?�����  ������Ĉ     |        A              >         �     Dp ����� ����� >�����  ����   � ?����� p   ��p     � ?����� }�               � ����� >�     8������� ?����� �?��������������� ����� A�����Ĉ     >        �                       A     Dq$���m�� ?����� }Ͷ�m�$�H�m�ܒI$�� ����� >�I$���x      � ����� ��               | ����� }�     x������� ��������������������� ����� �?�������            @              �        �      �x ����� ����� ������  ����   | ����� }�   �x|      | ���� �                > ����  ��     ��������� ���� ����������������� ���� ������     �       �              �       @    | ����| ���� �����  ����   > ����  ��   ��>      >  ��� �                  ?��� �     ���������  ��� ������������������ ?��� �������     �                      ��      �    >$���m�>  ��� �m�$�H�m�ܒI$�  ?��� �\�I$���        ��� �                � ��� �     ���������� ��� #�����������������@ ��� ��������    ��      "               �@            ����  ��� �����  ����   � ��� ��   ���     �  ��  �                �  �  �     ��������@  ��  G�����������������   �  #������$�@    �@      D                �       "     $������  ��  �����  ����   �  �  ��   ���     �      p                �      �     ��?������        ������������������      G������D�      �        �                |      D     Dč��m��      t���m�$�H�m�ܒI$���      �ܒI$����     �      >�                �      p     x�������      A�����������������       ���������     |      A                >       �      �������      >�����  ����   ��      w�   �x�     �      }�                 �      >�     >��������      �?�����������������      A�������     >      �                       A     A������      }�����  ����   ��      >��   �� �      �      ��                 |      }�     }��������     ������������������      �?�������          @                �      �      � ����m� �      �����m�$�H�m�ܒI$��|      }�ܒI$�}� |      |     �                  >      ��     �����������     �������������������     �������     �     �    ������     �     @     |���� |     � ����      �   �>      ���   �� >      >     �     ������           �     �����������     ������      ��������    ��������     �                �    ��    �     >���� >     � ����������x   �     ��   ��            �     �������     �    �     ������������    #������      ������@    ���������    ��    "           @    �@          ��m�$     �$���m���������I$���    �ܒI$��� �     �    �     �������     �    �     ����������@    G������      ?������     #������ ��@    �@    D                 �     "       ����� �    � �����������   ��    ���   �� �     �    p          �     �    �     ����?������      �������������������    G������@��      �      �      ������     |    D     @ ����� �    p ����     �   ���    ���   �� �     �    >�     >     �     �    p     ���������    A������������������     ����������     |    A     A������     >     �      � �I$�6��    >��rI$�>     �m��rI�    rI#m��_� �     �    }�     }      �      �    >�     >���������������?����������������������������� ��     >�����      �������     �����     A  �   ���    }���   }      �����  �    >� ������  �      �������     �      |      ������     }����������     �������������������    ?������ ��          @    �������     �          �   �   �����������   �      }����  ������ ���}��  |      �����     �      >      ?������     �������������    ��������������������    ����� ���     �    �    �������     �    @       |I$�6�`�����6�rI$��      >m��rI ?������I#m�����  >      ?�����     �            �����     �������������    ��������������������    ������ ���     �         ��������    �    �       >   ��?��������  �      ���  �����  ������                  �      �               ������������������������ ������������������������ ����    ������      �������@    ������           ��     ���  �      ����         ������  �               �      �               �����������������������@�������?�����������������  ���@    ������     @�������      ������         �$�6�l     ��rI$��      Ͷ�rI$     �I#m�����  �                     �               ������?������������������������������������������@ ���      ������      ��������     �����     @   �  ��     ���        ����         �����  �                >�      �                ���������������������� ������������������������� ���     �����     A �������     ?�����      �   �  ���    ���  >�      ����          �����  �                }�       �                >���������������������� ������������������������  ��     ?�����     � �������     �����     A    �$�6�m�    ��rI$}�       ���rI$�    �I#m�����   �                ��       |                }���?������������������ �������������������������  ?��                ��������                �     �  ���   ����  ��       }���   ���   ��}���   |               ��    �  >                ����������������������� �����������������������   ���                ��������                     |  ���   ���� ��       >���   ���   ������   >               ��   �                 ����������������������� �����������������������  @���                ���������                @   >$�6�m�$�I#m��rI#��       6�rI$�6�m�$�I#m�����                  ��   �  �              ��� �������������������  ����G������������������  �����                ��������@                �     ���   ���� ��  @  ���   ���   �����    �              ��   �  �              ��� ������������������@ ��������?���������������   ���@              @ ��������                     � ���   ���� ��  �  ���   ���   �����    �              �>  �  �              ��� ���?���������������� ����G������������������@  ���                � ��������              @     Ē6�m�$�I#m��rI� F  ��rI$�6�m�$�I#m����    �              >��  �  �              ��  ������������������  �����������������������   ���              A  ��������               �     � ���   ���� >��   ���   ���   ����    �              }���� �   �              >���  �����������������   ��������������������    ��              �  ��������              A      � ���   ���� }��    ���   ���   �����     �              �����  �   |              }���  ?����������������   ?���������������������    ?��              ���������              �       ��6�m�$�I#m��rH��� 
1   |�rI$�6�m�$�I#m}���     |             �����p     >              ����  �����������������  ?���������������������     ���              ���������                     | ���   �������"   >��   ���   �����     >             �����   �              ����  �����������������  ?��������������������  @  ���              ����������              @     > ���   �������<$  �   ���   �����                  ������׀� �            ���   �����������������    (h?���������������  �  ����              ���׀���@              �     6�m�$�I#m��rG������h  �rI$�6�m�$�I#k���      �            ������� ?� �            ���   ����������������@  (�����?�������������     ���@            @ ���� ?���                     ����   ������� ?����� ��   ���   ����      �            �����+ � �            ���   ���?��������������  ^4�����������������@    ���              � ��� ���            @       ����   ������ ���  ��   ���   ���      �            >���� p � �            ��    ����������������  �?t������������������     ���            A  �   }���             �       �6�m�$�I#m��r>������  �rI$�6�m�$�I#_��      �            }���>    �  �            >���    ���������������  �?8$�����������������      ��            �  >    |���            A        ����   ����}����?8��  ��   ���   ����       �            �����  �  x            =���    ?��������������  '�>8D�����������������      ?��              �  |���            B         ����   ���������>8D�� {�   ���   ����       |           ����� �  8            ;���    ���������������  w�L?������������������       ���             @�  ���            D          |6�m�$�I#m��q�����L8��� ;rI$�6�m�$�I#;���       >           ���  � ��  8            ;���    ���������������  ���������������������  @    ���             � `  ?����            D  @       >���   ���������p@   ;�   ���   ����                  ���  � ��  8            ;��     ���������������  �Q��������������������  �    ����               � ����            D  �       ���   ��������ќ��    ;�   ���   ���        �          ���  � ��  8            ;��     ��������������@ ���8�������������������      ���@          @    � �����            D         �$�H�m�ܒI$�������8���`  8���m�$�H�m�ܻ��        �          ���    p  8            ;��     ���?������������ ����?�����������������      ���            � �     q���            D         �  ����   ������9�  8����  ����;��        �          >����     �  8            ;��      ��������������  ��87 ����������������       ���          A  	�      ����            D         �  ����   >����`�87�  8����  ����;��        �          }���� ?�   <  8            ;��      �������������  ��0� ���������������       ��          �  �     <��            D         �$�H�m�ܒI$}���O�Dy0�<  8���m�$�H�m�ܻ��         �          ������?�    8            ;��      ?������������   ���� ?���������������       ?��           #� 
   ?��            D          �  ����   ����J��  8����  ����;��         |         ������?�  �  8            ;��      �������������  @����� ���������������        ���           C�    ���            D           |  ����  �����}��  8����  ����;��         >         �����   �  8            ;��      �������������  ������%?��������������� @      ���           ��@    ���            D @         >$�H�m�ܒI#����O����%?  8���m�$�H�m�ܻ��                  ��� �   �  8            ;�       �������������  �w��� ���������������� �      ����                 ���            D �           ����  �������"� 8����  ����;�          �        ��� �    À 8            ;�       ������������@  ?����e0���������������       ���@        @       Ã��            D          � ����  ���?���e3� 8����  ����;�          �        ��    8 �� 8            ;�       ���?����������  ?�����p|���������������       ���          �       ����            D          ĒH�m�ܒI��?�����p}� 8���m�$�H�m�ܻ�          �        >���    | � 8            ;�        ������������   �����x� ���������������        ���        A        ���            D          � ����  >��������x�� 8����  ����;�          �        }���8   8|   � 8            ;�        �����������  ������� ��������������        ��        �  8   8   ��            D          � ����  }���;�������� 8����  ����;�           �        ����8   ||  � 8            ;�        ?����������   ������ ?��������������        ?��          8   |   �?�            D           ��H�m�ܒH����;������� 8���m�$�H�m�ܻ�           |       ����p ��8  8p 8            ;�        �����������  @��}> � ��������������         ���         @p ��   8p�            D            | ���� ����q��} �p 8����  ����;�           >       ��� p �� �p 8            ;�        �����������  � ?��)���  ��������������@        ���         �p   �   p�            D@           > ���� ��� p>�)��< p 8����  ����;�                  ��� p �� � p 8            ;         �����������    ������ �������������Ā        �����������   p  �    p�            D�                  ��� p����p 8���m�$�H�m�ܻ            ����������� � �| � x 8   �����   :         ���        @   ������� �����    ����         ���        @  �  |  � x�   �����   E            ����������� �������x 8�����������:            ����������   �8 � 8 8     �    8         ���        � �?������� ����� � ����         ���        �    �8 � 8�   ��?��   F            �����������?�������8 8�����������8            ����������� � �  � 8 8     0    8          ���         ��������� ����� 0 ����          ���          � 	    � 8 �   �����   D            �������������������� 8���o�����m�ܸ                    ��� � �  �  8          8          ����������   ��������� G����   ����          ����������   �         D   �����   D                    ������<����� 8�����������8                    ��� � � �  8     @    8          ?����������    ��|����   G���� @ ����          ?����������    � �      D   �����   D                    ������|���> 8 8�����������8                    ����    :>   8     @    8          ����������  @ ������{�$ G���� @ ����          ����������  @ �    >   D   �����   D                    ����������{�< 8���o�����m�ܸ                    �� �     < 8     ��    8          ����������  � ��x�o� G���� �� ����          ����������  � �     8 D   �|}��   D                    �� ���h�o�< 8�����������8                    �� �8   �� < 8     ��    8          ����������   ��� N G���� �� ����          ����������   �8   �� 8 D   �x=��   D                    �� ���� N< 8�����������8                    �� �� �� < 8     �B    8          ����������   o���� G���� �B ����          ����������   �   �� 8 D   �x=��   D                    �� �o�<��� 8���o����m�ܸ                    �� � � �� > 8     ��    8          ����������   �����"  � G���� � ����          ����������   �    �� 8 D   ��=��   D                    �� �����"  � 8�����������8                    �� � � �� ~ 8     ��    8           ����������  ����   G���� � ����           ����������   �    �� x D   ��}��   D                    �� ��O�� ~ 8�����������8                    �� � �p�� v 8     @    8           ���������  �O����A� G����   ����           ���������   p  � �� x D   �����   D                    �� �O����]�~ 8���o�����m�ܸ                    �� ������ v 8          8           ?���������   �~���  � G���� @ ����           ?���������    p�  �� x D   �����   D                    �� �yO� �~ 8�����������8                    �� ������ v 8          8           ��������� @ �8��,"� G����   ����           ��������� @  p�  �� x D   �����   D                    �� �8'$"�~ 8�����������8                    �  ������ � 8      0    8           ��������� � �9��> @ G����   ����           ��������� �  8� P�� � D   �����   D                    �  �9<u" @� ;rI$�������I#8                    �  �� p�� � 8     �    8           ���������  �`?�|, p  G����   ����           ���������   8�   �� � D   �����   D                    �  �`?�,$ p � ;�  �����  �                    �  ��    � 8           8           ���������  �D?� �x  G����    ����           ���������   �    � D   �����   D                    �  �D?� �x!� ;�  �����  �                    �  �     > � 8           8           ���������  �;�� �� G����    ����           ���������        > � D           D                    �  �?�� ��� ;rI$�    �I#8                    �  �       � 8            8            ���������  �;��#��  G�������������            ���������          � D            D                    �  �;��#��� ;�   ���   �                    �  �       � 8            8            ��������  �#��#�   G�������������            ��������          � D            D                    �  �#��#� � ;�   ���   �                    �  ��      8            8            ?��������   ��� �  G�������������            ?��������    �      � D            D                    �  ���� o�� ;rI$�6�m�$�I#8                    �  ��       8            8            ��������@  ��(�  G�������������            ��������@   �      � D            D                    �  ���(�� ;�   ���   �                       �� �    8            8            ���������  �)��  G�������������            ���������   � �   � D            D                       ��)��� ;�   ���   �                        �� �   < 8            8            ��������   �  	#�  G�������������            ��������    � �   ?� D            D                        �� 	+�?� ;rI$�6�m�$�I#8                        �� �   � 8            8            ��������   �� 	7�  G�������������            ��������     x �   �� D            D                        �� 	7��� ;�   ���   �                        �� �  � 8            8                        �� 	7   G�������������                          | �  �� D            D                        �� 	7�� ;�   ���   �                         �� �  �8 8            8                         ��    8 G�������������                          > �  �� D            D                         ��  �� ;rI$�6�m�$�I#8                         �� �  �8 8            8                         ��    8 G�������������                           �  �� G�������������                         ��  �� 8            8                         ����   8 ?�������������                         ��    8 @                                      ��  �� @                                     ��� �� ?�������������                         ��    | p ?�������������                         �    p @                                      �    �� @                                     �� �� ?�������������                         ��    � � ?�������������                         �     � @                                      �    ��  @                                     ��  ��� ?�������������                         �~   � �                                        �      � �������������                          �   ��  �������������                         ��  ���                                        ?��   �                                        ?�      � �������������                          ��  ��  �������������                         ?���  ���                                        ?��  �                                        ?�     � �������������                           ��  ��  �������������                         ?���  ���                                        ?�����<�                                        ?��    <� �������������                           �����  �������������                         ?��������                                        �������                                        ��    �� �������������                          �����  �������������                         ���������                                        ������                                        �   �� �������������                           �����?�  �������������                         ���������                                        ���   �                                        ���   � �������������                           x�����  �������������                         ���������                                        ��� �                                          ��� �   �������������                           > ����  �������������                         ��������                                         ����� ?                                         ����� ?  �������������                           �  ��  �������������                         ��������                                         �� ��  ~                                         �� ��  ~  �������������                           � ���  �������������                         ��������                                         ��     �                                         ��     �  �������������                           �����   �������������                         ��������                                          ��    �                                          ��    �  �������������                           �����   �������������                          ��������                                          ��    �                                          ��    �  �������������                            �����   �������������                          ��������                                          ��   �    ���������                            ��   �  ��        ��                            ?����   ��        ��                          �������    ���������                            ?��   ?�    ���������                            ?��   ?�  ��        ��                            ����   ��        ��                          ?�������    ���������                            ��  ��    ���������                            ��  ��  ��        ��                            ���    ��        ��                          �������    ���������                            ��� �     ���������                            ��� �   ��        ��                             ��    ��        ��                          ������     ���������                            ��� ��     ���������                            ��� ��   ��        ��                             �     ��        ��                          ������     ���������                            ������     ���������                            ������   ��        ��                                    ��        ��                          ������     ���������                             �����     ���������                             �����   ��        ��                                    ��        ��                           �����     ���������                             ?�����     ���������                             ?�����   ��        ��                                    ��        ��                           ?�����     ���������                             �����     ���������                             �����             @                                                @                             �����     ���������                             ����      ���������                             ����              @                                                @                             ����      ���������                              ���      ���������                              ���              @                                                @                              ���      ���������                              ���      ���������                              ���              @                                                @                              ���      ���������                               ��       ���������                               ��               @                                                @                               ��       ���������                                        ���������                                                @                                                @                                        ���������                                        ���������                                                @                                                @                                        ���������                                        ���������                                                @                                                @                                        ���������                                        ���������                                                @                                                @                                        ���������                                        ���������                                                @                                                @                                        ���������                                        ���������                                                @                                                @                                        ���������                                                                                          ���������                                        ���������                                                                                                                                            ���������                                        ���������                                                                                                                                            ���������                                        ���������                                                                                                                                            ���������                                        ���������                                                                                                                                            ���������                                        ���������                                                                                                                                            ���������                                        ���������                                                                                                                                            ���������                                        ���������                                                                                                                                            ���������                                        ���������                                                                                                                                            ���������                                        ���������                                                                                                                                                                                                                                                             