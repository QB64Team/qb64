��`  |J� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         ����������������������������������������������������������������������������������������������������������������������������������������������������������������������� �                                       ������������������������������������������������������������������������������������������������������������������������������ ����������������������������������������������������������������������������������������������������������������������������������������������������������������������� �������������������������������������������                                       o���������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                               ����� p �������������������������������������������������������������������������������������������������������������������������������                               ����� p ����������������������������������    ����������������������������������������������������������������������������������������                               ����� p ����������������������������������    ����������������������������������������������������������������������������������������                               ����� p ����������������������������������    ����������������������������������������������������������������������������������������                            ����� p ����������������������������������    ����������������������������������������������������������������������������������������           p                ����� p ����������������������������������    ����������������������������������������������������������������������������������������           `                ����� p ����������������������������������    ����������������������������������������������������������������������������������������     8     8 �                ����� p ���������������������������������    �������������������������������������g����������������������������������������g�������� 8    0�    0�                 ����� p ��������������������������������    �������������������������������������'���������������������������������������'�������� 0    �    �                 ����� p ��������������������������������    �������������������������������������������������������������������������������������� 0   ��   ��                 ����� p �������� ?���� ?������������������    ��������������������������������������p������������ ?���� ?��������������������p������ `����!���� ?            ����� p ����>�|����|��~|���������������    ���������������������������������������&�������>�|����|��~|������������������&����� `����������ρ��           ����� p ����? ??�q�??�p>0~ ������������    �����������������������������������������������? ??�q�??�p>0~ ��������������������� �σ������c���           ����� p ���0|>?���>?��`�>������������    ���������������������������������������g�������0|>?���>?��`�>���������������g������ ��������8cw            ����� p ���>Dp�~�x��>�ǜ����������������    �������������������������������������$�&������>Dp�~�x��>�ǜ�����������������$�&����� ����1��pg�8?            ����� p ���<��|����|����������������    �������������������������������������fp�������<��|����|�����������������fp�������� 8`� `g�8            ����� p ���<������ǟ|��1���������������    �����������������������������������������������<������ǟ|��1����������������������������<x��ǌ             ����� p ���|9��������?8s���������������    �����������������������������������������������|9��������?8s����������������������������8�����            ����� p ���xq�����?���?0���������������    �����������������������������������������������xq�����?���?0������������������������� |<p�<�� �            ����� p ��������Ï����?1���������������    ����������������������������������������������������Ï����?1���������������������������p��9��8            ����� p ������q�����~a����������������    ��������������������������������������������������q�����~a����������������������������`;� �1��0�            ����� p �����y�?����?�|c� �������������������������������������������������������    ��������y�?����?�|c� ������������������������8���7��q�8q�                   p �����������xǎ��������������������������������������������������������������������������xǎ������������������������1� �<� a�0c�8                   p �����?���?�<����qϜ��������������������������������������������������������������������?���?�<����qϜ������������������������8q���x�� ��p��                   p ���ǎ��?�>���������������������������������������������������������������������ǎ��?�>��������������������������� �� �!�� @� A��                   p ����� ���~���߾ ?������������������������������������������������������������������� ���~���߾ ?�����������������������   �            �                    p ������������������ ��������������������������������������������������������������������������������� ������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������@  @  @      �       @         p ���������������������}����������������������������������������}�����������������������������������������}����������������������
@  @  @         �       @         p ���������������������}����������������������������������������}�����������������������������������������}�����������������������@  @  @         �       @         p ���u�����������������}����������������������u�����������������}�����������������������u�����������������}�����������������������X�OX�N
�����2�p��̐X����,r'  p ���t�����q��?q�?9���O�v3o��cwӍ�������t�����q��?q�?9���O�v3o��cwӍ��������t�����q��?q�?9���O�v3o��cwӍ�������JeQdQQ!Q �)J��"�"�(�e��2
(� p �����뮛���������uֵuw�7�u�o����]w����������뮛���������uֵuw�7�u�o����]w�����������뮛���������uֵuw�7�u�o����]w��������JEQDQ_j-_��$"��"�>S�E���"yO� p �����뮻��������u��u�w��o���]w݆��������뮻��������u��u�w��o���]w݆���������뮻��������u��u�w��o���]w݆�������EQDQP
!P@�"��"� R�E ��"�H  p ���5�뮻���������u��u�w߭�o����]w�v�������5�뮻���������u��u�w߭�o����]w�v��������5�뮻���������u��u�w߭�o����]w�v�������*E�DQQ
!Q �)J��"�""(`E"�"��� p ���պ�.����������uֵuw�w��ן�����g�ww�����պ�.����������uֵuw�w��ן�����g�ww������պ�.����������uֵuw�w��ן�����g�ww�����)D�ODNN
 �N���2�p�!�@D��h"x�  p ���ֻ����������?9���w��7����݇x������ֻ����������?9���w��7����݇x�������ֻ����������?9���w��7����݇x������               �         @         p ����������������������������������������������������������������������������������������������������������������������������               �        �          p �������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                         @       p �������������������������������������������������������������������������������������������������������������������������������  $                     @       p �������������������������������������������������������������������������������������������������������������������������������  $                     @       p ��������������������������������������������������������������������������������������������������������������������������������6s�9c��$q�+��6rG�"��IX��  p ����8Ɍ�iƜq�gێ0���ct�ɍ��8�L�1����cw�������8Ɍ�iƜq�gێ0���ct�ɍ��8�L�1����cw��������8Ɍ�iƜq�gێ0���ct�ɍ��8�L�1����cw������ �(��Y�QP(�(��������(��QId��  p ���}�[u���k����u�S]�]u�[uw}�]5������]w������}�[u���k����u�S]�]u�[uw}�]5������]w�������}�[u���k����u�S]�]u�[uw}�]5������]w�������/��=P0�訢��$����QUD��  p ���}�[��������W]�]u��t�}�]u������]w������}�[��������W]�]u��t�}�]u������]w�������}�[��������W]�]u��t�}�]u������]w�������($�EP(�����$����QUD��  p ���}��}�������}�W]�]u��uw��]u������]w������}��}�������}�W]�]u��uw��]u������]w�������}��}�������}�W]�]u��uw��]u������]w�������(��QEQP$�(��"���H�(��Q"D"�  p ���}�[u�������u�W]��e�[u�}�Yu��ݻ���g������}�[u�������u�W]��e�[u�}�Yu��ݻ���g�������}�[u�������u�W]��e�[u�}�Yu��ݻ���g��������r�=��"q�(�jr'���"Dh  p ���|8��n��q�oݎ0�a������8�v�1ݻ���������|8��n��q�oݎ0�a������8�v�1ݻ����������|8��n��q�oݎ0�a������8�v�1ݻ���������                                  p �������������������������������������������������������������������������������������������������������������������������������               <                   p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������      �              � �><� 
    p ����������������������������0�������������������������������������0��������������������������������������0������������     �              �$ �B�    p �����������������������������^�������������������������������������^��������������������������������������^�����������     �              �$ �@�    p �����������������������������^�������������������������������������^��������������������������������������^�����������<�8���r/��Ng fq�V�5��@�z��  p �����i�N?���O���ߙ���O�q��^��vg��������i�N?���O���ߙ���O�q��^��vg���������i�N?���O���ߙ���O�q��^��vg������ ��DY� �(��%Q@��
(�T�&Q��@���P  p ���]u���5�u�}7�뮿_k��[�7ٮ�oA��uu�������]u���5�u�}7�뮿_k��[�7ٮ�oA��uu��������]u���5�u�}7�뮿_k��[�7ٮ�oA��uu���������D����(���G�Dz/�T�$_�@���  p ���]u���t}�}w�`�_���o�w۠��^��uv�������]u���t}�}w�`�_���o�w۠��^��uv��������]u���t}�}w�`�_���o�w۠��^��uv���������E� �(��	�H�$�(T�$P�@�"���  p ���]u����u�}�}w��o�_�u���wۯ��^��uwo������]u����u�}�}w��o�_�u���wۯ��^��uwo�������]u����u�}�}w��o�_�u���wۯ��^��uwo��������EQ� �h��%H���(���$Q�B�"��P  p ���]u���u�u�}w���_ku�[�kwۮ��^��ue�������]u���u�u�}w���_ku�[�kwۮ��^��ue��������]u���u�u�}w���_ku�[�kwۮ��^��ue���������8���q���G�by���N!<�zi�  p ���C�n�v?�P�w��_����mw�����ᅖw������C�n�v?�P�w��_����mw�����ᅖw�������C�n�v?�P�w��_����mw�����ᅖw������  �                                 p ����������������������������������������������������������������������������������������������������������������������������  �               �                p ���������������������?���������������������������������������?����������������������������������������?���������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                    p �������������������������������������������������������������������������������������������������������������������������������   �    �                          p �������������������������������������������������������������������������������������������������������������������������   �    �                          p ��������������������������������������������������������������������������������������������������������������������������,��rH�Տ                         p ���8�?�����*p�����������������������������8�?�����*p������������������������������8�?�����*p�����������������������������	(�� ��H%�Q                         p ����M��}u���i�������������������������������M��}u���i��������������������������������M��}u���i������������������������������	/��������Q                         p ����]�}uW�k�������������������������������]�}uW�k��������������������������������]�}uW�k������������������������������	("����	�Q                         p �����~��}uW��k��������������������������������~��}uW��k���������������������������������~��}uW��k������������������������������	(����%�Q                         p ����]~��}v���k�������������������������������]~��}v���k��������������������������������]~��}v���k������������������������������	'"@��q�TO@                        p ����ݿ�}�����������������������������������ݿ�}������������������������������������ݿ�}����������������������������������                                     p �������������������������������������������������������������������������������������������������������������������������������                                     p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������O>��  �  ��        �     @  p �������{�����������������������������������{������������������������������������{�������������������������������P��$ H  @   $    � 	       p ���w������������������������������������w�������������������������������������w������������������������������������P��D$  H  @   $    � 	       p ���w�������������������������������������w��������������������������������������w�������������������������������������
P��D��c�� M��A�[fp5��`��+c��V8 p ����w}��J~�l~��cS������q�q�4���p��������w}��J~�l~��cS������q�q�4���p���������w}��J~�l~��cS������q�q�4���p�������
P��D�A�TA�I�AR��&QA@�,��	�AQYD p ����w��Y�k����M���kwٮ���u�S]�k�鮦�������w��Y�k����M���kwٮ���u�S]�k�鮦��������w��Y�k����M���kwٮ���u�S]�k�鮦������	P����AW�I�AR�$_@�訢	��QQ| p ����w�W[��>��]����w۠��tW]��>���������w�W[��>��]����w۠��tW]��>����������w�W[��>��]����w۠��tW]��>��������Ј���ATI"�AR�$P@���	QQ@ p ���/w�W[�����]����wۯ��u�W]������������/w�W[�����]����wۯ��u�W]�������������/w�W[�����]����wۯ��u�W]������������Ј��ATAI"�A��$QQ@�(��	AQQD p ���/w��[�뫾��]��-��wۮ���u�W]��뮮������/w��[�뫾��]��-��wۮ���u�W]��뮮�������/w��[�뫾��]��-��wۮ���u�W]��뮮������O��A���E�A�IpN�@�Ȩ���OQ9 p �������k��l��]������p�7Wa��������������k��l��]������p�7Wa���������������k��l��]������p�7Wa����������            @  A                     p �������������������������������������������������������������������������������������������������������������������������������               �                     p �����������������~����������������������������������������~�����������������������������������������~��������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������� �( @            @          p ����{���������������������������������������{����������������������������������������{��������������������������������������$  H            @       p ����������������������������������������������������������������������������������������������������������������������������D$   H            @       p ���������߷���������������������������������������߷����������������������������������������߷���������������������������������D��c�� O4�� 	9vD�Y���psN9����� s  p ����J~�l߰�1���3�c>S�ጱ�c>]M8ߌ�������J~�l߰�1���3�c>S�ጱ�c>]M8ߌ��������J~�l߰�1���3�c>S�ጱ�c>]M8ߌ������D�A�T@@H�Q 	EIE(e"�2�"�QE"�"�(�
  p ����Y�k����Z����ﶺ���~�w�u���~�4�_��������Y�k����Z����ﶺ���~�w�u���~�4�_���������Y�k����Z����ﶺ���~�w�u���~�4�_���������AW�@H�_ 	EID�E>�"�"�_A"�"�/�z  p ���W[��?��Z����ﶻw��~�����~�u�_�������W[��?��Z����ﶻw��~�����~�u�_��������W[��?��Z����ﶻw��~�����~�u�_���������AT �H�P 	EIDHE �"�"�PA"�"�( �  p ���W[����Z����ﶻ���~��}���~�u��u������W[����Z����ﶻ���~��}���~�u��u�������W[����Z����ﶻ���~��}���~�u��u�������AT@�H�Q E0IM(E"�"�"�QE"�&�(��  p ����[�뫿�Z����϶����~�w�u���~�u�_u�������[�뫿�Z����϶����~�w�u���~�u�_u��������[�뫿�Z����϶����~�w�u���~�u�_u�������A���O$��$8�I4�D���prN8����' y  p ����k��l��1���/��;�c]�፱�ceu�߆�������k��l��1���/��;�c]�፱�ceu�߆��������k��l��1���/��;�c]�፱�ceu�߆������        @  @(                        p �������������������������������������������������������������������������������������������������������������������������������          �@                        p ����������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������          !              �      p ����������������������������������������������������������������������������������������������������������������������������	    �    @!                   p ����������������������������������������������������������������������������������������������������������������������������	    �    @!                   p ����������������������������������������������������������������������������������������������������������������������������c������c�`!98���Y��89��9����   p ���~XS>'�i������?N3�So���'�~4�N8�������~XS>'�i������?N3�So���'�~4�N8��������~XS>'�i������?N3�So���'�~4�N8�������	�A(��%�Y@?ED �(e)�%E,��(�  p ���k��M~��k��������5����o�������}5�������k��M~��k��������5����o�������}5��������k��M~��k��������5����o�������}5�������	�(��%��@!E|��(E)��<=%�E���  p ����>�]~��h.�޺���u���o�������au��������>�]~��h.�޺���u���o�������au���������>�]~��h.�޺���u���o�������au�������	(��%�@!E@@�(E)�DE% E��   p ������]~��k�޺����u����o�������]u�����������]~��k�޺����u����o�������]u������������]~��k�޺����u����o�������]u��������	A(��%�Q@!ED �(E)`DE%E(��(�  p �����]~��k��޺����u���럻�����]u���������]~��k��޺����u���럻�����]u����������]~��k��޺����u���럻�����]u��������'�A$䓑(!98���D��@<=$�9Ȟ��   p ����~�]��ln������?v;�W�������7av8��������~�]��ln������?v;�W�������7av8���������~�]��ln������?v;�W�������7av8�������    �                  @             p ����������������������������������������������������������������������������������������������������������������������������                     �             p ����������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                     @     @�   p �����������������������������������������������������������������������������������������������������������������������������            ��       � `0  �  0 p ���������������?�������?�����<�������������������������������������������������������������������?�������?�����<�������������            �       � @` �    p ����������������������������{��������������������������������������������������������������������������������{�������������            �      � �@ ��  ` p �����������������������g�3���w��w������������������������������������������������������������������������g�3���w��w����������                   ��� � 0 @ p �������������������������?�����g��������������������������������������������������������������������������?�����g����������    �   `#�@ � ��`	0p�#8� p �������������������{��x��s��������<���������������������������������������������������������������{��x��s��������<�������   �   �i�6L�� ��  3�gd�0 p ����������������_�ɳ?�=���b_�������r������������^�����������������������������������������������_�ɳ?�=���b_�������r�������        |� hI�� {  `/ ^��  p ����������������4�����9������������{f������������������������������������������������������������4�����9������������{f�������cG�     �@xY�� �@@@{ ���  p ����������������i���{���!�������zM������c����}�������������������������������������������������i���{���!�������zM������"�����    u��[ 1�`3��@Fr �.` p �����������������?�/���{���j?��﹍��џ������k}wm�8�������������������������������������������������?�/���{���j?��﹍��џ������B� �   p� �� c�c? @0�f �x@ p ����������������0��h���?�������3��1������]���m��_�����������������������������������������������0��h���?�������3��1�������!� �  � � c �, @`���`  p ������������������@�����y���O;�u�������]��w���_�������������������������������������������������@�����y���O;�u����������H��   :8��: � h�@����2F  p �����������������?�\��9�����?��?3�e͹������]k}�s��^������������������������������������������������?�\��9�����?��?3�e͹������c'��  �i�9�v � i�!���fL� p ���������������=��Y��e������~>s�噳?���������|�����������������������������������������������=��Y��e������~>s�噳?�����           �� 1d � N ���p� p ���������������q����	��������~w��;������������������������������������������������������������q����	��������~w��;������     0                               p �������������������������������������������������������������������������������������������������������������������������������                                     p �������������������������������������������������������������������������������������������������������������������������������                                     p �������������������������������������������������������������������������������������������������������������������������������                                     p �������������������������������������������������������������������������������������������������������������������������������                                     p �������������������������������������������������������������������������������������������������������������������������������                                     p �������������������������������������������������������������������������������������������������������������������������������                                     p �������������������������������������������������������������������������������������������������������������������������������                                     p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p ���������������������������������������������������������������������������������������������������������������������������������������������������������������������� ��                                      ?����������������������������������������������������������������������������������������������������������������������������� ����������������������������������������������������������������������������������������������������������������������������������������������������������������������� �������������������������������������������                                       ��������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         ������������������������������������������������������������������������������������������������������������������������������