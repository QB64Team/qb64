�'k  �0� }                                                                                                                                                                                                                                   8                        8                                                 x                                                ~                        `                        �                        �                       ��                                               �                      ��                       �                      �                       ��                      �x                      ��                       a�                      ��                      �                      ��                       `                      ��                      ��                     ���                                           ��                     ���                     ��                      �                      ���                     ��x                     ���                       a�                     ���                     ��                     ���                       `                     ���                     ���                    ����                                           >��                    '����                    ?���                     a�                     ?���                    y��x                    ?���                    F  a�                    � g�                    ~� �                    � g�                    a `                    e� �                    | �                   g� ��                   �                     � �                   � ��                   � �                   H �                    � ��                   � �x                   � ��                    H  a�                   z  g�                   �  �                   �  g�                    $  `                    z  �                    �  �                   �  ��                   $                      =  �                   o  ��                   }  �                     �                    =  ��                   o  �x                   }  ��                      a�                   �  g�                   7�  �                   >�  g�                   	   `                   �  �                   7�  �                  >�  ��                  	                      @  �                  �  ��                  @  �                  �  �                   @  ��                  �  �x                  @  ��                  �   a�                  �  ��                  ������                  ������                  @   `                  �����                  ������                 ������                 @  �                  �����                 �  ���                 �����                 �����                  ���� ��                 ������x                 ���� ��                    �a�                 ���� '�                 ������                 ���� '�                  �  ��`                 �    �                 ������                �    ��                 ������                  ������                 ��������                �������                 @    �                  �    ��                �    �x                �    ��                 H     a�                 z     g�                 �     �                 �     g�                 $     `                 z     �                 �     �                �     ��                $                      =                      o     ��                }     �                     �                 =     �                o     �x                }     ��                     a�                �    '�                7�    ��                >�    ��                	     `                �     ��                7�    �               >�    ���               	     �                @     ��               �    w��               @    ��               �     ��                @    A��               �    ��x               @    ��               �     Pa�               �     @G�               �    ���               �     �g�               @    @�`               �     �)�               �     ���              �     �y��              @     (�               �      &�              �     ����              �     pv�                    ���               �     PA��              �     m��x              �     x��                    Pa�              �     @g�              x     m��              �     8�g�               �     UP`              �     ��              x     7`�             �     =���              �     
�               �     (��             �     7`��             �     ?��              H     ��               �      ��             �     ��x             �     ���              H     @ a�              z       g�              �     � �              �     � g�              $     @ `              z     
  �              �     � �             �       ��             $     �               =        �             o     � ��             }       �                  � �              =        ��             o        �x             }        ��                      a�             �        g�             7�        �             >�        g�             	         `             �        �             7�        �            >�        ��            	                      @        �            �        ��            @        �            �        �             @        ��            �        �x            @        ��            �         a�            �         g�            �         �            �         g�            @         `            �         �            �         �           �         ��           @                     �         �           �         ��           �         �                     �            �         ��           �         �x           �         ��                      a�           �          g�           x          �           �          g�            �          `           �          �           x          �          �          ��           �                      �          �          �          ��          �          �           H          �            �          ��          �          �x          �          ��           H           a�           z           g�           �           �           �           g�           $           `           z           �           �           �          �           ��          $                      =           o�          o           ��          }           �                     �           =           ��          o           ��          }           ��                      @           �           ?�          7�           �          >�           �          	                        �           ?�          7�           ��         >�           ��         	                       @           ?�         �           ��         @           ��         �                      @           ?��         �           �x         @           ��         �            �         �           ?��         �           ���         �           ���         @            `         �           _��         �           ���        �           ����        @                     �           o��        �           ����        �           ���                     �         �           ���        �          ���x        �          ����                      a�        �           � g�        x          � �        �          � g�         �             `        �           � �        x          � �       �          � ��        �                      �          � �       �          � ��       �          � �        H             �         �          � ��       �          � �x       �          � ��        H              a�        z          �  g�        �          �  �        �          �  g�        $              `        z          �  �        �          �  �       �          �  ��       $                      =          �  �       o          �  ��       }          �  �                     �        =          �  ��       o          �  �x       }          �  ��                      a�       �         �   g�       7�         �   �       >�         �   g�       	               `       �              �       7�         �   �      >�         �   ��      	                      @          @   �      �         �   ��      @         `   �      �              �       @              ��      �         �   �x      @            ��      �               a�      �               g�      �         ,h    �      �         #�    g�      @               `      �         �    �      �         ;�    �     �         $H    ��     @                     �         �    �     �         ;�    �      �         $H    �                     ��     �         �          �         ;�    ��     �         $H    ��                             �                �     x         ,h     �p     �         #�     ��      �                      �                �     x         �     �     �              ��      �                �      �               �     �         �     �     �         `     ��      H                �      �                �     �         �    �     �         �    ��      H                �      B         �    �      �         �    ?�p      �         �    ?��                                      �    ?       �         �   ���      �         �   ���                              !         �   �        _         �   ���      m         �   ��                     8�                 �   �                �   ~?�       N         �   �       1              ��                 �   ��       �        �  ���                �  ���        �                      �        �  ��        �        �  ��        �        �  ��         @             p8         @        �  �8        �        �  ��        q�        �  ��8                     ��                  �  ���        �        � ���        n�        � ���                                      � ��         {�        � ?�         Up        � ?��         *�            �p                 � ?�p         q�        ����         _h        ���p          �           �                 ���         {�        ����         Ud        ���         *�           8                 �|�          �    ����~?�          .�    ����          Q        ��           �    �� ���          �   ?��������          1��   ?��������          N	                      /P   ?� ���           ?��   ?� ����           �p   ?� ����            �         p8           ��|   |  �~8           �������������           �߃���������8           S          �            ����������q�            ?�����������            ������������            (�                      	����������             �|   |  ��             	�����������             �������� p             ?���������p             �����������             ?����������             �                        ǃ���������             �����������              �����������             8                        8        |               ?���������               8        �               ��������                ���������               ���������               ���������                                        ��   �                  ����                   �    �                                           �������                        �                  ������@                                           ~    �                        @                  ~    �                                                 �                                                 �                                                 `                                                 `                                   