��g  X  ��������������������������������������p��p��p��p��p��p��p��p������������� �� �� �� ����������������������������������������������������������?��?��?��?��?��?��?��?���������������������������������������������������������                                                                         /  .  �   � X� ?    \  ^  9    �  �  v  0  j b  �  ` p x  �  ` � � �  � � � � � � � � � � � `   �   �     � @   /@ .@ �   � X� ?    \  ^  9      9        
                                                 y          