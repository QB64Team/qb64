�h  �z��                 `                                              `                                              `                                              `                                             �` 0                                           �` 0                                           �` 0                                           �` 0                                            ` 0                                            ` 0                                            ` 0                                            ` 0                                           g�8<��ny����<��<                               g�8<��ny����<��<                               g�8<��ny����<��<                               g�8<��ny����<��<                               3lٰf��l��m���f                               3lٰf��l��m���f                               3lٰf��l��m���f                               3lٰf��l��m���f                               �o�0f�������0>͛~                               �o�0f�������0>͛~                               �o�0f�������0>͛~                               �o�0f�������0>͛~                                                                                                                                       �l03f�����͛0f͛`                                                                                                                                                                                           �lٰ3f́�l͛m�0f͛f                                                                                                                                                                                           g�<���fy���0>��<�                                                                                                                                                                                                                                                                                                                                                                                                                           �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ?��                ��                ��                                                                                                                                                                       � |                �               | �                                                                                                                                                                      x  �             �                �  <                                                                                                                                                                     �   8                 �             8   �                                                                                                                                                                                     0                 �    `                                                                                                                                                                    0    �            �                                                                                                                                                                                         �     `                �                                                                                                                                                                                                          `           0     �                                                                                                                                                                                   0                 �      `                                                                                                                                                                                   @                                                                                                                                                                                                 �          �                                                                                                                                                                                         �       `                �                                                                                                                                                                                                          @                                                                                                                                                                                                                             �                                                                                                                                                                                                  @        @                                                                                                                                                                                                   �                                                                                                                                                                                          @                                                                                                                                                                                                   �        �                                                                                                                                                                                         @         @                                                                                                                                                                                                 �                           �                                                                                                                                                                                                          @                                                                                                                                                                                                                             �                                                                                                                                                                                                           �                                                                                                                                                                                              @          @                                                                                                                                   @                                                           �                                                                                           @                                                  �                                         @                                                                                                           �                                                  �                                         @                                                                                                           �                                                                                      �      �                                                                                                                                                                                                �      �                                                                                                                                                                                    @           @                                                                                                                                                                                     @     @           @                                                                                                                                   @                                                 �     �                             �                                                                                                                  �                                                       �                             �                                                                                                                                                                                                      @                                                                                                                               @                                                                       @                                                                             @                                                  @                                                                                          �                                                            @                                                  �                  @                                                                       �                                                            �                  @                               �                  �                                                                        �                                                            �                  �                                                  �                  @                                       @            @                                                                              �                  @                                                 �                                       @            @                                                                                                �                                                                                        @            @                                                                                                                                                                                        @            @                                                                                                                                                                                         �                                                                                                                                                                                           �          �                                       @                                                  �                                                 H                  �            `                 �          �      �             0                  �                  �             X                  x                               P                 �                 `            l                x          �     �             x                 �                 �                               �                  `             �                  �                 �            �                ~          �                  �                 �                 �             (                 �                  �             �                                  �            �          @     �               8            �                                  �             (                 �                 �            D                                  �           �          @     �               x           �                                  �             P                 �                 �            D                                   @           �          @     �               �           �                                  �             P                 �                              �                                  .�           �         @     �               1�           ��                ?                 ?�             �                 �                 @            ��                                 ]<           �         @     ��              c��          ��                �                �            �                 �                 �            �                �                ��          �?�        @     7���             ǃ�          ���               o��               ���           G�                /�                 9|            ��               ?��              t��          ���        @     /��            ���         ���               0���              ����          @>                 �                r�           
'��               `_��              ���         ���       @     _��?�           ���         g���              q����             ���          ��               . �               �           
8?��                ���             Ӄ��         ����       @     �����           ?���        x?��              a����             �����         ��               �_ <              �| �          W���              @���             �|��        ����      @     ����?�          ���        �����             �����            �|��          > �              | ��             ��          `~��            ���?��            N���        ����      @    �����          ����       �~��            ǁ�?��            �����        �              �@�<             )  �         (����             �����            ����       7����     @    ���~          �����       =�����           �����            ����        
  �            �@ <�            I  �         (� ��           � <?�            @ ���       7� ���     @    �� ?���         �� ��?       =� ��           � <?��           _@ ���        
H  �            �  �p            �� �        Q�  ���           � ���           @ �       o�  ��~     @    �� ���         �� ���      {�  ���           � ���           �@ ��       H  �           �   <            �  �8        z  �            �  <�            �  ���      �  ���     @     �x  ?�?         �  ���      �  ��           �  <�           �  ���       $   �p            �  ��           "@          z   ���           ��  ��           @�  ?�      ^   ���           yx  ���     �     �  �       z   ���           9�  ���           �  ?�       $               ��   p8           @@  ��       =   �          �   q��          ��  ��       o   �>           �   ��     �     �  ���       }   �           �   q��           �  ���         ��           H              �    8        =   ��           �   ?�          �   8��      o   ��           �   �8     �     �   ?��       }   ��           �   ?�           �   8��           p0           H   ��                      �   q�           z   ��          �   �      7�   �            �   ��     �     x   �        >�   q�            �   ��           �   �       	               $    80           �    ��      @�   <           z    8�          �    ��      7�   �            �    ?�     �     x    ��       >�   <            �    8�           �    ��      @	    �           $                �           @@   �           =                �    �      �   �           o    �     @     �    �       @   �            }                �    �      @�    0                �           H           �@    0           =     �           �           �    <           o     �     @     �    �       @    0            }     �           �           ��                                H     �      ��               �                 z     �      �               7�    0     @      �     �       �                >�                 �     �      �@                	                  $            �                 �              @  z            �               7�         @      �     @       �                 >�                 �            @                 	               @  $            �                 @              �  =            �               �                 o     �       �                 @                 }                              �              �              �               @ @                =            �               �                 o     �       �                 @                 }                            @ �                            �               � �                �           x               �                 7�    �       �                 �                 >�            �               � @                	            �               � �                �           x               �    @           7�           �                 �                 >�            �               � @                	             �                �                @           �               �    @           �           �                 �                 @            H                                 �            �                �                @      �     �                �    �           �           �                 �                 @            H                                 �            z                �                 �      �      �                x    �           �            �                 �                 �            $                 �                 @            z                �             @   �      @      �    @           x               �            �                 �                 �            $                 �             @   @            =                 �             �   �      @      o    @           �               �            }                 �                 �                             H             �                 =                 �                �             o    �      �     �               �            }                 �                 �                              H                              �                z                �             7�   �      �      �               x            >�                 �                 �             	                 $                 �          @  �                 z                �            7�         @      �               x            >�                 �                 �          @  	                  $                 �          @  @                 =                 �            �         @      o               �            @                 }                 �          @  �                                  H          �  @             @   =                 �            �                o          �     �             @                 }                 �          �  �             @                    H          �  �             �   �                 z            �               7�         @      �   @         �                 >�                 �          �  @             �   	                  $            �             �   �           @     z            �               7�                 �   �         �                 >�                 �            @             �   	            @     $            �                @           �     =            �               �                 o   �         �                 @                 }                             �           �                 �                @                =            �               �  @             o            �                 @                 }                             �                            �                �                �      �     x                �  �             7�           �                 �                 >�            �                @                	            �                �                 �      @     x  @             �               7�           �                 �                 >�            �                @                 	             �                �                 @            �  �        �     �               �           �                 �                 @            H                                  �            �                �                 @           �          @     �               �           �                 �                 @            H                                  �            z                �                 �            �                x          �     �             �                 �                 �            $                 �                 @            z                 �                 �            �               x          @     � @           �                 �                 �            $                  �                 @            =                  �                 �            o               �                 � �           }                 �                 �                              H                               =            @     �                 �            o               � @              �            }                 �                 �                         @     H                               �           �     z                 �       �     7�`               ��              x            >�                 �                 �             	            �     $                  �        @    �                 z                 �             7��          �     �               x            >�                 �                 �        @    	                  $                  �        @    @                 =                  �            �           @     o               �            @                 }                 �        @    �                                   H        �    @                 =                  �            �           0     o           �    �`            @                 }                 �        �    �                                   H        �    �                 �                 z            �                7�           0     ߀            �                 >�                 �        �    @                 	                  $             �                                   x        �    �                7�                �             �                 >                  �                                                                                                            0    �            �                     x                                                 `                                                                                                                                 0                 �    `                                                                                                                                                                    �   8                 �             8   �                                                                                                                                                                     x  �             �                �  <                                                                                                                                                                      � |                �               | �                                                                                                                                                                       ?��                ��                ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      � `�  ��         ̀`             �         0                                                                                                                                                              0    ��         l `�             0     0                                                                                                                                                                 0    ��          `�             0     0                                                                                                                                                                 1�n�><��;`<��<     �|�y�<��y�      ��͹��3π                                                                                                                                                            1��lٻ�����f     ͳv�Ͷf���      ͳ3m�m�7m�n�                                                                                                                                                            1��lٳ>����>͛~      m�f���~��͘      3?m��3�f6l�                                                                                                                                                            1��lٳf����f͛`      m�f���`�f͘      30m�3c6l�                                                                                                                                                            1��lٳf���`f͛f     m�f�ͶfͶ͘      �3m�m�6m�l�                                                                                                                                                            1��f�3>��30>��<     ͟f`y�<��y�      �m�͙�g3��                                                                                                                                                                                                                                                                                                                                                                                      �        >                                                                                 