�i  l�g�                             �       `�  l                                                            �       `�  l                                                            �       `�  l                                                            �       `�  l                                                            0       ��  l                                                            0       ��  l                                                            0       ��  l                                                            0       ��  l                                                                    ��  l                                                                    ��  l                                                                    ��  l                                                                    ��  l                                                            ������p<��������p                                                         ������p<��������p                                                         ������p<��������p                                                         ������p<��������p                                                         �m�6 `�`f���m�0l�                                                         �m�6 `�`f���m�0l�                                                         �m�6 `�`f���m�0l�                                                         �m�6 `�`f���m�0l�                                                          7�����`f���6m�3�`                                                          7�����`f���6m�3�`                                                          7�����`f���6m�3�`                                                          7�����`f���6m�3�`                                                                                                                                                                                                                    6�`͛`f�͛6m�6l0                                                                                                                                                                                                                                                                                                6m�6`͛`f�͛6m�6l�                                                                                                                                                                                                                                                                                                �������`<���3����sl                                                                                                                                                                                                                                                                                                      �                                                                                                                                                                                                                                                                                                                   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                          �                 �                 (        @        
         P        �                 �                 (        @        
         P                                                                                                                                                                  �                 �                 (        @        
         P        �                 �                 (        @        
         P                                                                                                                                                                  �                 �                 (        @        
         P        �                 �                 (        @        
         P                                                                                                                                                                  �                 �                 (        @        
         P        �                 �                 (        @        
         P                                                                                                                                                                  �                 �                 (        @        
         P        �                 �                 (        @        
         P                                                                                                                                                                  �                 �           �     (        @        
         P        �                 �           �     (        @        
         P                                                                                                                                                                 �                 �          ?�     (        @        
         P        �                 �          ?�     (        @        
         P                                       �                                                                           �                                            �                 �           �     (        @        
         P        �                 �           �     (        @        
         P                                       �                                                                            �                                            �                 �           �     (        @        
         P        �                 �          �     (        @        
         P                                        x                                                                                                                         �                 �           p     (        @        
         P        �                 �          p     (        @        
         P                                                                                                                                                                �                 �           8     (        @        
         P        �                 �          8     (        @        
         P                                                                                                                                                                �                 �                (        @        
         P        �                 �               (        @        
         P                                                                                                                                                                �                 �                (        @        
         P        �                 �           �     (        @        
         P                                        �                                                                                                                       �                 �                (        @        
         P        �                 �           G     (        @        
         P                                        �                                                                                                                       �                 �           �    (        @        
         P        �                 �           #�    (        @        
         P                                         �                                                                            �                                           �                 �           8    (        @        
         P        �                 �           8    (        @        
         P                                         �                                                                            8                                           �                 �           �    (        @      
         P        �                 �           �    (        @      
         P                                        �                �                                                         �                                           �                 �           �    (        @ �     
         P        �                 �           �    (        @ �     
         P                                        �                �                                                         �                �                         �                 �           �    (        @      
         P        �                 �           �    (        @ /     
         P                                         �                ��                                                         �                                         �                 �           �`   (        @      
         P        �                 �           �   (        @ ]�     
         P                                         q                >�                                                         `                                         �                 �           ��   (        @ �    
         P        �                 �           �    (        @ ��    
         P                                                         x �                                                                           �                        �                 �            ��   (        @ ��    
       P        �                 �            �    (        @ ��    
       P                                         0@               p p        �                                                0                  @                        �                 �            s�   (        @ P �    
  �     P        �                 �            x   (        @P �    
  �     P                                         0�               � 8       ��                                               0                @         �               �                 �            �   (        @` p    
  �     P        �                 �               (        @p p    
  �     P                                         1�               �        ��                                                               @        �               �                 �            3�   (        @� 8    
  ��    P        �                 �            0   (        @��8    
  .�    P                                         @               �        �                                                               �         �              �                 �            |   (        @ �     
  
�    P        �           �    �               (        @ �8    
  K�    P                                                        �        < p                                                               �         @              �            @    �            >   (        @ @     
  T �    P        �            `    �  �           (        @ �    
  T �    P                     �                                  �      8 8                                                                                        �           �    �              (        @ �     
  ( p    P        �           �    �           �  (        @��    
  � p    P                     �       �                        � �      p                            �                                  �                        �           0`    �  �        ��  (        @ � �   
  � 8    P        �           0`    �  �        �@  (        @� C�   
  � 8    P                     ��       �                       �  �      `                            0`       �                         �  �                      � ��        PP    �           �  (        @ � �   
  �     P       ���        ]�    �            `  (        @� �   
  ��    P  00      >         �<       �         �             �  p      `        �                  @                                 �  @      @               ���        �8    �  

        �x  (        @ �  �   
  @     P  ?�    ����       �8    �  �        ��  (        @� 0�   
  ~    P  ��     ��        �       <�         �x             �  8      � �      �      ��         �                 �               �         @        ?�     � `      �    �           ��  (        @ �  p   
    �   P  x0    � x      �    �           �   (        @� p   
  p�   P x0     ���               p�         ��             �        � �      ��                                 �               �           �      x0     �a��      �    �  8�        ��  (        @ �  8   
  ` �   P  �(    �,��      �    �  8�        �   (        @�  8   
  � ��   P ��     ��        �      � �        ��             �        @ �     �       �                 �         �               �        @ �      �     � =           �  p�       �p  (        @ �     
  ` �   P  �    �[ ?=�          �  p�       �   (        @�    
 p >x   P �     <  �        �     � p        �p             �        � �     �        <               @ @        �               �        @ x      �     �t  g@      �   �  � �       @   (        @ �     
  ` �   P @    �t �`     |�   �  � �       @   (        @�    
 p �   P @     8  �      8  �     � 8         �              �  �     � �     ��     0           �      �                           �        @ �           �(  �      �   � � p            (        @ �  �  
  ` ��  P �    ��  =�     ���   � ��p            (        @ �  �  
 p �   P 
�     p  �      p  p                               �  �     � �      �        �        @                                �   �     @ �           �0  t       �   � � 8            (        @ �  �  
  ` ��  P  �   ��  v     8 `�   � �p8            (        @ �  ��  
 p �   P ��    `   �      �  |                               �  �     �  @       �         p                                         �  �     @          �    ��   ]     0  �   �   �           (       @ �  �  
  ` �@  P  �   ����݀    � �   �  �           (  ��   `@ �  .x  
 p ��  P >�    `   >        �       �                      �  �     �  �       p     @            �       �                        �  x     @  �       @    ��   @    � �   �    �           (    ���@ �  �  
  ` π  P   �   �� ?�w`   � �   �  ?�           (  �� @@ �  �  
 p �@  P ���    @   �    �  �        �                 ���  �  �     �  �       8     @         �  �        �                 �     �  �     @  �            ��   	�   � ��  �    ?�  ����������    � 0@ �  �� 
  `  O�  P    N   ��  <�   � ��  �    ��  ����������   }���@@�  �  
 p  `   P  0N        �       �       �             ����� 0  �  �     �  �       >         �       w�       �                 �     �  �     @  @            �`   O   � �0  �    ?�           �������@ �  �� 
  `  ��  P      ��  O   � �@  �    >�           ����� @@@�  �  
 p  �  P  �    @   ��   
   8�       �             �������  �   @     �  e            @    G       0        �             �����     �         @  @           ��   �     ��  �    ?�  �����������������@ �  �@ 
  `  e�  P   ��  ��   �?�     �   �    >�  ��������������� @@@�  �� 
 p  `  P  �   @    ��                               ���  �   �     �  0�      �    @    �                                 �     �   �     @          g�   ��    ��     �  �    �           (����ß�@ �  π 
  `  0�  P   ��  ��   0��     ~  �    �           (������ @@�  �@ 
 p  0  P '  ��   @    ;�   0                              �  �   �     �  @      ?�    @    3�                                         �   �     @         ;�   ��    ��     9�  �    �           (    ��0@ �   �� 
  `  |  P   ��  ��   ��     <  �    �           (    �� @@�   �  
 p    P '  ��   @    ��   `   @                         �0  �   �     �         @    @    ��                                  �    �   �     @             ��    ��  (   	�  �    >           (     �@ �   �� 
  `  >  P   �  ��   ��  �     �    �           (     <s�@@�   � 
 p    P   {�   @    �   `   �                        �   �   e     �             @    ?�                                       �   `     @              �@    ��� P   �  �    ?           (      @@ �   u� 
  `   @ P   ?�  ��    �  �     �    ��          (      `@@�   p 
 p   � P   ?        y�      �                           �  �   0�    �  @                                                   @   �   0     @              �     z~` �   �  �    ?�          (       �@ �   8� 
  `  � P   �  �     {�� `     �     @          (       �@ �   8 
 p    P           ~`             �                    �  �   @    �  �                                                     �   �        @             �     ��       �    ��          (        @ �   | 
  `  � P    �  �     �`      � �    �           (       �@ �    
 p     P           �              �                    @  �        �  �     `                           �                        �        @              �     �     � �     ��          (        @ �   > 
  `  � P    �  �            @ �     �          (        @ �    
 p     P            ��      �        a                       �       �  �      P                          @                        �        @              �     ��     �� �     a�          (        @ �   @
  `  � P    _  �           �  �     `          (        @ �   �
 p     P     �       ���      �        0�                      �   @   �  �                        �                                 �        @              �     ���      � �     8�          (        @ �   �
  `     P    � �     �       0 �     8          (        @�    
 p     P     @       ���      �       @                      �   �   �          �         �                                         �        @               �      �w�      �� �      y          (        @ �   �
  `      P    �� �     �      �@ �                (        @�     
 p      P    �         `w�      @�       !                      �   �   �            �          `        @                                 �        @            �   �      p?�      @� �     7�         (        @ �   �
  `      P     �� �      p       @  �               (        @�     
 p      P     �        0?       @|       �                     �   �   �            A          0        @                                �        @            @   �      8      @| �     �  0      (        @ �   �
  `      P     � �      x       @  �         |      (        @�     
  p      P                     �|       �                     �   �   �            `�                 @                                �        @                �      (       �8 �     �  A�     (        @ �     
  `      P     `� �      (       �  �         A�     (        @�     
  p      P     `                 �8       �   >                 �        �             ^                 �                                �        @                �             �  �        �     (        @ �      
  @      P      ~ �      8       �  �         �     (        @�      
  �      P                       @            �                �                       >                               �                 �                          �                �         |9    (        @ �      
         P      > �                �         X|9�   (        @�      
         P                                     '��               �                      p>                                 |                �                          �                �          #��    (        @ �      
         P     ` �                �          ��    (        @ �      
         P     `                                 ?��              �                      p                                 �                �                      `   �                �           �   (        @ �      
         P     P  �                �          q�w�   (        @ �      
         P     P                                  ��              �                                                           g�               �                          �                 �            �a�  (        @ �      
         P        �                 �          �   (        @�      
         P                                         ���                                                                          �                                           �                 �           �~  (        @        
         P        �                 �           ����� (        @        
         P                                        �x                                                                         �                                           �                 �            ��� (        @        
         P        �                 �              (        @        
         P                                        ���                                                                                                                     �                 �            r��� (        @        
         P        �                 �           �   (        @        
         P                                         ��                                                                                                                     �                 �            �� (        @        
         P        �                 �            ;@  (        @        
         P                                         ��                                                                                                                     �                 �            �� (        @        
         P        �                 �            �   (        @        
         P                                         �                                                                           �                                          �                 �             �� (        @        
         P        �                 �            �   (        @        
         P                                          p                                                                                                                      �                 �             (   (        @        
         P        �                 �             l   (        @        
         P                                                                                                                                                                �                 �                (        @        
         P        �                 �                (        @        
         P                                                                                                                                                                �                 �                (        @        
         P        �                 �                (        @        
         P                                                                                                                                                                �                 �                (        @        
         P        �                 �                (        @        
         P                                                                                                                                                                �                 �                 (        @        
         P        �                 �                (        @        
         P                                                                                                                                                                 �                 �                 (        @        
         P        �                 �                 (        @        
         P                                                                                                                                                                  �                 �                 (        @        
         P        �                 �                 (        @        
         P                                                                                                                                                                  �                 �                 (        @        
         P        �                 �                 (        @        
         P                                                                                                                                                                  �                 �                 (        @        
         P        �                 �                 (        @        
         P                                                                                                                                                                  �                 �                 (        @        
         P        �                 �                 (        @        
         P                                                                                                                                                                  �                 �                 (        @        
         P        �                 �                 (        @        
         P                                                                                                                                                                  �                 �                 (        @        
         P        �                 �                 (        @        
         P                                                                                                                                                                  �                 �                 (        @        
         P        �                 �                 (        @        
         P                                                                                                                                                                  �                 �                 (        @        
         P        �                 �                 (        @        
         P                                                                                                                                                                  �                 �                 (        @        
         P        �                 �                 (        @        
         P                                                                                                                                                                  ��������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           ?����������                                                                  ?����������                                                                  ?����������                                                                  ?����������                                                                                                                                                                                                                            ?����������                                                                                                                                                                                                                                                                                                         ?����������                                                                                                                                                                                                                                                                         �     @  � ��   @            ?����������  
      @  @     
�  P �                                                                                                                                                                                                                                             P       � ��  �@         ?����������  
      �  @      �  @ �                                                                                                                                                                                                                                                   � ��  �@         ?����������       �  @      �  @@                                                                                                                                                                                                                                            䁬p"sND�������N03��A�s��  ?����a���� �,�����Ec��x�'"
��S�C�9�                                                                                                                                                                                                                                          2�"
QE �,���(�QH$A"A2�H"�  ?��ݺ뮿��� (���� �E�@D(�
� TT$QE                                                                                                                                                                                                                                          "�zQD��袾���_ $A"A"�H"�  ?��ݾ�.���� 
�/���S��E@�D�(�
��T$}                                                                                                                                                                                                                                          "��QD@�(���(�P$A"A"�H"�  ?��������� 
�("��R �EAE(�
� T�A                                                                                                                                                                                                                                          U�"��QM �(���(�QH$A!�"�H"�  ?����뮿��� B(�"�" �MAE Ȧ
� TRQE                                                                                                                                                                                                                                          ��@�pzN4��螜��DN0�� �rHi  ?����a���� B'"h!��5��x� �
��S��9�                                                                                                                                                                                                                                                                        ?����������              @  �                                                                                                                                                                                                                                                                                  ?����������              @                                                                                                                                                                                                                                                                                       ?����������                                                                                                                                                                                                                                                                                                         ?����������                                                                                                                                               ?����������                                                                  ?����������                                                                                                                                                                                           