��a  \m�            �0     `   �     � �                       �0     `   �     � �                       �0     `   �     � �                       �0     `   �     � �                       �0        �    � �                       �0        �    � �                       �0        �    � �                       �0        �    � �                        0        �    � �                        0        �    � �                        0        �    � �                        0        �    � �                       3ǜ�o��l�fx���<�8                      3ǜ�o��l�fx���<�8                      3ǜ�o��l�fx���<�8                      3ǜ�o��l�fx���<�8                      ��l��6m�ll�f��6c3fٰ                      ��l��6m�ll�f��6c3fٰ                      ��l��6m�ll�f��6c3fٰ                      ��l��6m�ll�f��6c3fٰ                       ߷��6m��l�<��7�0fٰ                       ߷��6m��l�<��7�0fٰ                       ߷��6m��l�<��7�0fٰ                       ߷��6m��l�<��7�0fٰ                                                                                                                   �6�6m�ll�<��60fٰ                                                                                                                                                                ٶl��6m�l8��s6l3fٰ                                                                                                                                                                �3ǌ��m��0�xc��<�0                                                                                                                                                                          0     c                                                                                                                                                                                �    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             ��                                           ��                                                                                                                                       ��                       ?�          ��     ��          ��                      ��     ��          ��                      ��      ��                                   ��                 @          �          ��     w           ��                      ��     ��          ��                    ��                                          ��               ��          ��          ��               P                    P     ���          ��          8          ��                  @                    P   ?�            @          ��          ��   �?�           ��                      ��   ����          ��                    ��    ?�                                     ��  8����         �           ��          �� ������         ���                      ��  ��� c         ���                    ���   ���                                     �� 1�����         ��         ���         �� �������         ����                     �� �����c         ����        �          ���� �����                                   ������o�        x��        ����        � �����o��       ����                    � � ������        ����       ����        ���� ���o�                                 � ����l       ���       �����       � �����|�      �����          |        � ��������       �����      ����       ������??�`          �           |        � ������}t�     ����      ?�����     �� ���7����}|�    ������         �      ��  ��??��߃�     �������      0?����     �������??��p          �          �      ��  ��/������X�    ������     �������      ����/������\�    ��� }�         ��        }|������|�     �������     �����     ������������|X          }|          ��        }|�����{��     �������    3�������      ����`_���?���@   ?�� ���         ��         ��`?����}�{�   ?�������    �������    ?���������?y�8          ��          ��         ��`������@   ?�������    �������    ���� ��`�������@   �� ��?�     >   ��    ��   �>`7����w���   ��������    #�������    ��������7����w��     �   �>      >   ��    ��   �>`?����G��@   p�����    � ����    ��  � ��������@   
� ��  �                
�       o���G��   ��������    w�������    ��������/���G��                            
�       ���^���    c�����    �>?���    ��    �������    ������          �     �    � o�������   �������    '������    �������o�����                             �       g���?���    �����  @    |���     �      ��������   ����<x`         ǀ         <x ���?��    �����Ç�    �����8|    �����Ç�G��>��                                     ���`�m��   �������    ?�����|~    <��Ǡ���������   ����?��    >`  7��    3�  �����      �����`    ����� $    �����`���                                         _� ��   ��������    >?���|~    a�
���Ǡ?���>����   ���|����    �� +��    � �����  �
 �    � ����`     ��� t    � ����`     
 �        ��                  �� ` ����   ��������    >>?���|~    c����Ǡ&���H�\!�   ���}���    ��p7��    �����  ���    � ����`     ��� $    � ����`              �          p         �   }�3�z�=�   ��������    >>?���|~    c�
���Ǡ@�]�~�_��   ���|����    �� ?��    � ������3�:�2    � ���@@    8 ���D    � ���@@              �                      �   ��H��<���   �������    8���8    ���`�����o]�   ����>p�    ��  �     �   p`�' D��    �#���㏀    >"?���8�    �#���㏀      @           `                         �����/���   � ���  �    8"���           `���������   ������    ��   �        �` D T b    �������    >>?����    �������      @           `                         �x���р   �����      <���     �     ��z������   �9�����     �   |     8   �� ��  * �    ������?     ?�����    ������?       �           �                         _�����+     ������     ?�������    8   ����������+�   ��������    ��  ��    ?�   ��� A
  5��     ������     ?�������     ������      �     8   ���    ��  ��     8   �� G�������    |�����     ��������   �   ���������π   �������    ��  ��    ��   }�>  }0    |�����     ��������   |�����       |     �   }�    ��  ��        }| #�� �    ������p    ���������   ��������{�� 1�   
��   ��     ��  �    
��   �� T��`    ������p    ���������   ������p  @         
��   ��     ��  �    �   �  ���x <    ?������     ���������   ��������|���x<?    ��   ��     >    |     ��   ��������    ?������     ���������   ?������  ��x       ��   ��     >    |      �   � 0~          �����      s�������         �p:~   ~    ?������p                     �p�������     �����      s�������     �����   .               �p                            p     �����      �������         � �� �     ������                      � ����      �����      �������     �����                   �                          LSU��                  �����      ������ �7�����     ������                  ������ �@(                     �����                           ������                          ޣ �                                       ޣ ��                                       �!\��                                                                                       }����^                                        �����_�                                       �����                                        ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    0 � 0`      �0 `�       �        �0 `�                                                                                                                                            1�   0       �6 `        �`        �6 `                                                                                                                                             00   0       �6 `        �`        �6 `                                                                                                                                             0><��l�     �7�ٞ      ��p>��     �7�ٞ                                                                                                                                           0;݃6lـ    ��lٳ      ��`f͛0     ��lٳ                                                                                                                                           03>ك6g��    ߶l�?      ��`f���     ߶l�?                                                                                                                                           03fك6g�     �6l�0      ̓`f��      �6l�0                                                                                                                                           1�fك6c�    ٶl�3      ͛`f�c0     ٶl�3                                                                                                                                           3>ف�c     �3��      ��0>�a�     �3��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �     �       >          �          �                                                                                                                                               P     �       !          (          P                                                                                                                                                    �       !          (                                                                                                                                                         g;,�       !9Y�        )�$        g;                                                                                                                                            H����       >e         �(�        H��                                                                                                                                            H����        =E         )�0        H��                                                                                                                                            H����        EE         *((        H��                                                                                                                                            QH����        EE         *(�        QH��                                                                                                                                            �G$�"�        =D�        ��"        �G$�                                                                                                                                                                                                                                                                                                                                          0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                < �     @ p�     � �                                                                                                                                                          "�      @ �$    � @                                                                                                                                                          "�      @ $    � @                                                                                                                                                          "r���pr'39NI�s9f��@                                                                                                                                                          <����"�(��EQI0"��E����@                                                              ���                         ����            ���                         ����                "���� �O�EQU"��}"��@                                                                                                                                                              "���� �H!EQU"��A"��@                                                                                                                                                              "����"����EQ"�"��E���@                                                                                                                                                              <r@�pp�#9N"p�r9��@                                                                                                                                                                                      @                                                                                                                                                                                      �                                                  