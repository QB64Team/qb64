��c  �-�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   P                                                                     P                                                                     0                                                                                                                                          �                                                                     �                                                                     p                                                                     0                                                                    `                                                                    `                                                                     �                                                                     `                                                                    �                                                                    �                                                                    �                                                                     �                                                                    �                                                                    �                                                                    �                                                                    �                                                                    `                                                                    p                                                                    �                                                                                                                                         �                                                                    �                                                                                                                                                                                                              -�                                                                    -�                                                                                                                                                                                                              [@                                                                    [�                                                                    <                                                                                                                                          ��                                                                    ��                                                                    x                                                                     0                                                                    m                                                                    o                                                                     �                                                                     `                                                                    �                                                                    �                                                                    �                                                                     �                         �      �    0    �                        �                        �      �    0    �                        �                        �      �    0    �                        �                         �      �    0    �                        �                        3 � `    �       �                        h                        3 � `    �       �                        x                        3 � `    �       �                        �                       3 � `    �       �                                                 0 � `    �       �                        �P                       0 � `    �       �                        �P                       0 � `    �       �                         0                       0 � `    �       �                                                0<�p<�6��3�7ǀ�6�                        -��                       0<�p<�6��3�7ǀ�6�                        -�                       0<�p<�6��3�7ǀ�6�                         p                       0<�p<�6��3�7ǀ�6�                         0                       fٳ`���6��l��6ـ                       [A`                       fٳ`���6��l��6ـ                       [�`                       fٳ`���6��l��6ـ                       < �                       fٳ`���6��l��6ـ                        `                       ~߰`>����3�o��6߀                       ���                       ~߰`>����3�o��6߀                       ���                       ~߰`>����3�o��6߀                       x�                       ~߰`>����3�o��6߀                       0 �                                                                  m�                                                                  o�                       `�0`f�͛1��l f6�                        ��                                                                   `�                                                                  �`                                                                  �p                       3fٳ`f��͛v��l��ـ                      ��                                                                   �                                                                   ��                                                                  ��                       <�0>�6���7ǀ��6�                     �                                                                   �                                                                   h-�                                                                  x-�                                                               �                                                                                                                                       �[@                                                                  �[�                                       p                         <                                                                                                                                       -���                                                                  -ව                                                                   x                                                                    0                                                                   [Am                                                                   [�o                                                                   < �                                                                    `                                                                   ���                                                                   ���                                                                   x�                                                                   0 �                                                                  m�                                                                  o�                                                                   ��                                                                   `�                                                                  �h                                                                  �x                                                                  ��                                                                   �                                                                   ��                                                                  ��                                                                  �                                                                   �                                                                   h-�                                                                  x-�                                                                  �                                                                                                                                       �[@                                                                  �[�                                                                   <                                                                                                                                       -���                                                                  -ව                                                                   x                                                                    0                                                                   [Am                                                                   [�o                                                                   < �                                                                    `                                                                   ���                                                                   ���                                                                   x�                                                                   0 �                                                                  m�                                                                  o�                                                                   ��                                                                   `�                                                                  �h                                                                  �x                                                                  ��                                                                   �                                                                   ��                                                                  ��                                                                  �                                                                   �                                                                   h-�                                                                  x-�                                                                  �                                                                                                                                       �[@                                                                  �[�                                                                   <                                                                                                                                       -���                                                                  -ව                                                                   x                                                                    0                                                                   [Am                                                                   [�o                                                                   < �                                                                    `                                                                   ���                                                                   ���                                                                   x�                                                                   0 �                                                                  m�                                                                  o�                                                                   ��                                                                   `�                                                                  �h                                                                  �x                                                                  ��                                                                   �                                                                   ��                                                                  ��                                                                  �                                                                   �                                                                   h-�                                                                  x-�                                                                  �                                                                                                                                       �[@                                                                  �[�                                                                   <                                                                                                                                       -���                                                                  -ව                                                                   x                                                                    0                                                                   [Am                                                                   [�o                                                                   < �                                                                    `                                                                   ���                                                                   ���                                                                   x�                                                                   0 �                                                                  m�                                                            o�                                                             ��                                                                   `�                                                            �h          �                      �                 �        �x                                                            ��                                                             �                                                             ��          @                      @                 @        ��          �                      �                 �        �                                                             �           �                      �                 �        h-�    .      �                .      �           .      �        x-�    �     �                �     �           �     �        �           �                      �                 �                    �                      �                 �        �[@    ]�     �                ]�     �           ]�     �        �[�    >      �                >      �           >      �         <           �                      �                 �              Z�     
�                Z�     
�           Z�     
�        -���    Z�     �                Z�     �           Z�     �        -ව    =      �                =      �           =      �         x            �                       �                  �         0     1      `                1      `           1      `        [Am     ��     h                ��     h           ��     h        [�o     |      �                |      �           |      �        < �     0       `                0       `           0       `         `     0       h                0       h           0       h        ���     �      h                �      h           �      h        ���     z      �                z      �           z      �        x�     0       `                0       `           0       `        0 �     �      0                �      0           �      0       m�     �      �                �      �           �      �       o�     x      x                x      x           x      x        ��     `       0                `       0           `       0        `�     h       4                h       4           h       4       �h     j      �                j      �           j      �       �x     �      x                �      x           �      x       ��     `       0                `       0           `       0        �      `                      `                 `             ��     j      Z                j      Z           j      Z       ��     �       �                �       �           �       �       �      `                       `                  `              �      `                       `                  `              h-�     h      Z                h      Z           h      Z       x-�     �       �                �       �           �       �       �      `                       `                  `                             �                        �                   �       �[@     *       �                *       �           *       �       �[�     �       ^                �       ^           �       ^        <                                                                       (                       (                  (              -���     *       �                *       �           *       �       -ව     �       ^                �       ^           �       ^        x                                                                 0      �       F                �       F           �       F       [Am      �       V�               �       V�          �       V�      [�o      |       /                |       /           |       /       < �                                                                 `              �                       �                  �      ���      �       V�               �       V�          �       V�      ���      ~       /                ~       /           ~       /       x�                                                                0 �      !       #                !       #           !       #      m�      ��      +@               ��      +@          ��      +@     o�      ^       �               ^       �          ^       �      ��                                                                `�      J�      @               J�      @          J�      @     �h      Z�      +@               Z�      +@          Z�      +@     �x      '       �               '       �          '       �     ��                                                             �       ��������               ��������          ��������     ��      ]��������               ]��������          ]��������     ��      #�      �               #�      �          #�      �     �       �      �               �      �          �      �     �       `     �        �     `     �          `     �     h-�      .`     �        �     .`     �          .`     �     x-�      ��������         @     ��������          ��������     �        `      �                `      �           `      �             �������        <(     �������          �������     �[@      ������
�        �(     ������
�          ������
�     �[�      ��������        �     ��������          ��������      <        ������ �                ������ �           ������ �              �      �       ��      �      �           �      �     -���      �     ��       ��     �     ��          �     ��     -ව      ?�������        ?�     ?�������          ?�������      x               �        �             �                  �      0       ?������`       �?�     ?������`          ?������`     [Am       �������Eh      �?�     �������Eh          �������Eh     [�o             ��       ��           ��                ��     < �               `        ?�             `                  `      `             �h      �           �h                �h     ���       ?������h      ?�     ?������h          ?������h     ���        �     ��       ���      �     ��           �     ��     x�              �`       �            �`                 �`     0 �        '�������0     ���      '�������0           '�������0    m�        �������Ҵ     ���      �������Ҵ           �������Ҵ    o�             3�x      ���           3�x                3�x     ��              �0       ��            �0                 �0     `�              �4     �`            �4                 �4    �h              zҴ     ~��            zҴ                 zҴ    �x              �x     ���            �x                 �x    ��               �0      �               �0                  �0     �               a    �� �            a                 a    ��              aR    ���            aR                 aR    ��              �     ��@            �                 �    �                `     �                `                  `    �               `    <�h            `                 `    h-�              i[    |�x            i[                 i[    x-�              �    �����            �                 �    �                `     � @             `                  `                     h	   ����`             h	                  h	    �[@              h��  ����x            h��                h��   �[�              �^    ?����            �^                 �^     <                `    �  �@             `                  `                    0�  8?�<�0            0�                0�   -���              ���  �?���p            ���                ���   -ව              xN   �����            xN                 xN     x                0    ?� �              0                  0     0                4N� ����               4N�                 4N�   [Am               �^� ���� `            �^�                �^�   ��o               x'   ��?���            x'                 x'    < �                0   � �               0                  0     `               � ��x?� �            �                �  ���               Z]����?� �            Z]�                Z]�  ���                �#� �����              �#�                 �#�   x�                �  � ?�               �                 �   0 �                g����               g�����            g���m�               Z.g���� �            Z.g�����           Z.g���o�                �� ������              ��                 ��  ��                 ` � �                 `                  `   `�                � �����              �                 �  �h                � ������             �                 �  �x                ^�������               ^������            ^������                  �� �                                     �                  ���� p                ������             ����t�                ����?� ��             �������            �����|�                ^?�������               ^?�����            ^?����                  �� �                  �����             ���                  F� ��� �             F�                 F�  �-�                V�� ������             V��                 V��  �-�                /�����                /�����            /���                       ��                                                           ������              �������            �������@                V��������              V�������            V��������                / @ ���                 / @                 / @    <                     �                                                            #@0�� p�               #@0                 #@0   r�                +@���� ��               +@������            +@�����s�                � ?���                 �                 �    �                    �                                            p                 	���?��                	�������            	�������                 -���?���                -�������            -�������                 � ���                  �                  �    �                 �  ?�                   �                  �    �                 � ���                 �                  �    
                 � ����                �                  �                     	�����                   	������             	�������                  � �                     �                   �                      ���@?                  �����             �����4                 �����                 �����             �����<                 �����                   ������             �������                  ���                     �����              �����                     �                                           �                 �  ��                  �                  �     �                 ?���                    ?�����             ?�����                                                                                        ����                   ������             ������`                 �����                   ������             �������                                                                                                                                                          x �                    x                  x    �                 ���                    �����             ������                  �                        �                   �                                                                                              ?��                      ?�����              ?�����                   ����                     ������              ������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                0   `                � 0  0               � �                                                                                                                                                                                                                                    0   `                �                   l3 �                                                                                                                                                                                                                                    p   `                                   l0 �                                                                                                                                                                                                                                    s��>|y��             �3�7ǀ             l�0<���                                                                                                                                                                                                                                   �l��v��0             ���n��l�             m�f�6                                                                                                                                                                                                                                   ��ϳf͛�              ُ�l��o�             m�`͛6                                                                                                                                                                                                                                   �ٳf͛               ٙ�l��l              m�`͛6                                                                                                                                                                                                                                   �lٳf͛0             ٙ�l��l�             m�3f͛6                                                                                                                                                                                                                                   3�Ͼfy��             �����7ǀ             ��<���                                                                                                                                                                                                                                      �0                     `                                                                                                                                                                                                                                                             �0                    �                                                                                                         