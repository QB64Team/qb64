�n]  Ta�                                                                         ������������������������������������                                                                                                            ������������������������������������                                    ������������������������������������                                    ������������������������������������                                    ������������������������������������                                    ������������������������������������                                     ?����������                   ���� ��         ?�������������������   � ?����������                   ����                                     ������������������������������������                                    ������������������������������������                                     ?����������                   ���� ��0       ?�������������������   � ?����������                   ����   0                                ������������������������������������  0 0  �                        pp  ������������������������������������  0 0  �                             ?����������                   ���� ��0 0  �   ?������������������� 8�� ?����������                   ���   0 0  �                            ������������������������������������  7�;�<���                     �  ���������������������������������?��  7�;�<���                          ?����������                   ���� ��7m�3f͛��?������������������� �� ?����������                   ���   7m�3f͛��                         ��ə�̟2d���������������������������                                   ������������������������������������                                     ?ɜ�̟2d��                   ���� ��         ?������������������� �� ?����������                   ���                                     ��ɒLș2d�?�������������������������                                �  ���������������������������������?��                                     ?ɘ��Ó��                   ���� ��         ?������������������� 8�� ?����������                   ���                                     ������������������������������������                                pp  ������������������������������������                                     ?����������                   ���� ��         ?�������������������   � ?����������                   ����                                     ������������������������������������                                    ������������������������������������                                     ?����������                   ���� ��         ?�������������������   � ?����������                   ����                                     ������������������������������������                                    ������������������������������������                                    ������������������������������������                                    ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                      �(     P                                                      ������������������������������������                                      �(  $    �    �     @                                              ������������������������������������                                      DH  $    �    �     @                                              ������������������������������������                                      DK�5����Փ,q��NE��i��4�r                                        ������������������������������������                                      DL��&QU �T�� �QEAJP(�@�                                        ������������������������������������                                      *���$_V��R"� �QEI�%@�                                        ������������������������������������                                      *���$PU@�Q"� �QE �H�(%@�                                        ������������������������������������                                      ��$QT� �T�� ��MQJR(�@�`                                       ������������������������������������                                      ��N�N��S"q�N5�)���Hq�                                       ������������������������������������                                                                                                         ������������������������������������                                                                 0                                         ������������������������������������                                                                                                            ������������������������������������                                      �             @ @   �                                           ������������������������������������                                      �  	            @ @                                               ������������������������������������                                      �  	            "  @                                               ������������������������������������                                      �Ȝc��r�s��5c��"%c�I0<�c��                                        ������������������������������������                                      �(�	�AR� �R ��@"%�QIH"��QP                                        ������������������������������������                                      ��>	�R� ��@�EQU "���P                                        ������������������������������������                                      �% 	R� ��AEQU"��QP                                        ������������������������������������                                      �""	AR� �R(�A�Q"H"��QP                                        ������������������������������������                                      ����r r�Ǖ����"0<����                                        ������������������������������������                                                     @                                                    ������������������������������������                                                    �                                                    ������������������������������������                                                                                                            ������������������������������������                                            @ 
 �                                                     ������������������������������������                                              �                                                      ������������������������������������                                                                                                    ������������������������������������                                      IȰ9�sNX+rI������9c�`                                       ������������������������������������                                      J(�E"
Qd,��JA$��AYQQE�Q�                                       ������������������������������������                                      J(�A>zQD�(���$���_Q}�                                       ������������������������������������                                      J(�A �QD�(����$���QPQA                                       ������������������������������������                                      2)�E"�QDD(��A$��AQQQEQ                                       ������������������������������������                                      !Ơ9yNDD(�q�䤞�����9�                                       ������������������������������������                                                       �                                                  ������������������������������������                                      �                �                                                  ������������������������������������                                                                                                            ������������������������������������                                        �  �     �   @  �                                            ������������������������������������                                         @         @                                               ������������������������������������                                         @         @                                               ������������������������������������                                      rĂ�g		��y�8朰3�4[X��s��0                                        ������������������������������������                                      $��QH��+(ED��$P$Re	��J,�                                        ������������������������������������                                      z$�QH��(E@���$P$RE�	���K�                                        ������������������������������������                                      �$�QH�*(EA��$P$RE	��J�                                        ������������������������������������                                      �#QH�*(EE��$P$�E	��J(�                                        ������������������������������������                                      z"N'!�$y�8�#�#QD��rIȐ                                        ������������������������������������                                                A                                                          ������������������������������������                                                A                                                          ������������������������������������                                                                                                            ������������������������������������                                                    �                                                   ������������������������������������                                                    �	    �                                              ������������������������������������                                                    �	    �                                              ������������������������������������                                      s�X8r�0��r�͜r��,�����                                        ������������������������������������                                      �AdD�(H�"�
�)�)(��"
J)�                                        ������������������������������������                                      �D|�( �>�z���)/��"
J)�                                        ������������������������������������                                      �D@�("� ���)"�)("�"
J)                                        ������������������������������������                                      �QDD�(H"�"���)"�)(��"
J)�                                        ������������������������������������                                      r�D8r$0��z��r)'"@�
K��                                        ������������������������������������                                                                                                           ������������������������������������                                                                                                           ������������������������������������                                                                                                            ������������������������������������                                         !  @�                                                              ������������������������������������                                         @  @@                                                              ������������������������������������                                         @  @@                                                              ������������������������������������                                      IȰm9c�@                                                              ������������������������������������                                      J(�IE�R@                                                              ������������������������������������                                      J(�I}H@                                                              ������������������������������������                                      J(�IAD@                                                              ������������������������������������                                      2)�IER@                                                              ������������������������������������                                      !ƠI9�P                                                              ������������������������������������                                             @                                                              ������������������������������������                                      �      �                                                              ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                      �           � �  �   @                                          ������������������������������������                                                � @   �  �                                           ������������������������������������                                                � @   �  �"                                           ������������������������������������                                      !�s8�p-���$Y��1 g�"V<�                                        ������������������������������������                                      " �D��$@"���*(� H��"YE��                                       ������������������������������������                                      " �|���$�@ �0+�" O��TQER                                        ������������������������������������                                      " �A�"�%@ �(*" H"�TQEQ                                        ������������������������������������                                      " �E�"�%@"��*(�!H�� �QE$�                                       ������������������������������������                                      !�r8�p%$���"��GN �Q<�#                                        ������������������������������������                                                                                                         ������������������������������������                                                                                                          ������������������������������������                                                                                                            ������������������������������������                                      �     A       @�      �                                            ������������������������������������                                      ��    A      A                                                  ������������������������������������                                      ��     A      A                                                  ������������������������������������                                      �ݎxC��A��s�������X�c�(����                                       ������������������������������������                                      �AD �Q�AA�J)A"�d�A(�)�                                       ������������������������������������                                      ��OD �QUA��J)�A"��D���(�)�                                       ������������������������������������                                      ��QD �QUA�J)A"�E�(�)                                       ������������������������������������                                      ��QD �S%AA�J)A"�E�A)�)�                                       ������������������������������������                                      �ROy ��%A��rK�����D���&����                                       ������������������������������������                                         @                                                              ������������������������������������                                         @                   �                                           ������������������������������������                                                                                                            ������������������������������������                                      �      �  �   @      @                                         ������������������������������������                                      �           @      @                                         ������������������������������������                                      �           @      @                                         ������������������������������������                                      ����<�c�,p<�c��@�Y��4㔐x�                                        ������������������������������������                                      �)	EU�H2�"��Q�@R) �T�E                                        ������������������������������������                                      �)�	E��"�"���U@�R)'�ԐE�                                        ������������������������������������                                      �)	E"�"��QUAR)(�T�E                                         ������������������������������������                                      �)	EUH"�"��Q%A�)(�T`E                                        ������������������������������������                                      �$��<��"p<���%@�I�'���@x�                                        ������������������������������������                                                               @                                          ������������������������������������                                                              �                                          ������������������������������������                                                                                                            ������������������������������������                                           A      �@                                                      ������������������������������������                                         @@      �                                                       ������������������������������������                                         @@      �                                                       ������������������������������������                                      c�8�gY0<�=��Y�3�                                                   ������������������������������������                                      �QEH�eH"�E�$R(�Q                                                   ������������������������������������                                      C�}H�E "�E�S�$Q         �                                        �����������������������������������                              �      $JAH�E"�E"�R$Q     �   �                                        ��������������������������?��������                          �   �      �DEH�EH"�E"�$R(�P�   �   �                                        ����������������������������������                         �   �      c�8�'E0<�=�Q���   � � �                                        ��������������������������?�������                         � � �                        �    � �                                        ����������������������������������                          � �                x           �`fc                                         ���������������������������g��������                         �`fc                              wx��s                                         ��������������������������8������                         wx��s                              ����c                                         ��������������������������81������                         ����c                              ?����                                         ���������������������������33�����                         ?����                              <wq���                                         �������������������������È�# �����                         <wq���                              9�m���                                         ��������������������������9�b`8�����                         9�m���                              o�ǀ                                        ���������������������������`�8����                         o�ǀ                                1�                                         ������������������������������|�����                            1�                                 �                                         �����������������������������������                            �                                                                           ������������������������������������                                                                                                         ������������������������������������                                                                                                           ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                    