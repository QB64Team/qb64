�'k  �0� }                                                                                                                                                                                                          `                        `                                                                         �                        �                        f                        `                        ~                        �                        �                                              ��                       �                       `                                              ��                      ��                      �                       �                      ��                      g�                      �f                        `                      �~                      ��                       `�                                             ���                     ��                      `                                             ���                     ���                      �                       �                     ���                     �g�                     �f                        `                     9��~                     9���                     & `�                                            >ǟ�                    >��                    � `                                           ���                    ���                    ` �                      �                    �\ y�                    �| g�                    �  f                       `                    x� ~                    d� �                    �  �                    �                      � ��                   � �                   @  `                    @                      � ��                   � ��                   @  �                    @  �                   v  y�                   z  g�                    �   f                        `                    v  ~                    z  �                    �   �                                           ;  ��                   =  �                   P   `                                          ;  ��                   =  ��                   P   �                      �                   �  y�                   �  g�                   (    f                       `                   �  ~                   �  �                   (    �                                         �  ��                  @  �                      `                                         �  ��                  @  ��                      �                      �                  `   y�                  �  ��                  
��� f                       `                  ����~                  �����                  
     �                                        �������                 �����                 ��� `                 ���                   �������                 ���� ��                      �                      �                 �  ���                 ���� '�                 �     f                  �     `                 ������~                 �    �                 �     �                 �                       ���� ��                 �������                @     `                 @                       �    ��                 �    ��                @     �                 @     �                 v     y�                 z     g�                 �      f                        `                 v     ~                 z     �                 �      �                                        ;     ��                =     �                P      `                                       ;     ��                =     ��                P      �                      �                �    y�                �    g�                (     �f                      `                �    ~                �    9�                (     ��                                     �    ���               @    ��                    �`                     �                �    ���               @    ���                    ��                     ��               `     �y�               �    Pg�               
      ��f                     @ `               `     �>~               �    @�               
      �P�                    @               �     `7��              �     ���                    pp`                                     �     `1��              �     �)��                    x��                      �              �     0`y�              �     UPg�              �     8� f               �     @ `              �     0`~              �     PP�              �     =� �              �     @                �     ���              �     *��             @     � `              @     �                �     ���              �     (���             @     � �              @     � �              v     � y�              z     @ g�              �     �  f                       `              v     � ~              z     @ �              �     �  �                                    ;       ��             =     
� �             P        `                                   ;       ��             =     � ��             P        �                      �             �        y�             �       g�             (          f                       `             �        ~             �        �             (          �                                   �        ��            @        �                      `                                   �        ��            @        ��                      �                      �            `         y�            �         g�            
           f                       `            `         ~            �         �            
           �                                  �         ��           �         �                      `                                  �         ��           �         ��                      �                      �           �          y�           �          g�           �           f            �           `           �          ~           �          �           �           �           �                       �          ��           �          �          @           `           @                       �          ��           �          ��          @           �           @           �           v           y�           z           g�           �            f                        `           v           p           z           ��          �                                               ;           ��          =           p@          P            �                                  ;           ��          =           �           P            �                                  �           ?�          �           @          (            ?�                                  �           ?�          �           @          (            ?�                                �           ?�         @           @�                     ?�`                                �           ?��         @           @�                     ?�                      �         `           ?��         �           ��         
            ?�f                       `         `           _�~         �           �9�         
            _��                               �           o���        �           �F�                    o�`                               �           ���        �          ���                    � �                      �        �           � y�        �           g�        �           �  f         �              `        �           � ~        �           �        �           �  �        �                       �          � ��        �           �       @          �  `        @                       �          � ��        �           ��       @          �  �        @              �        v          �  y�        z            g�        �          �   f                        `        v          �  ~        z            �        �          �   �                               ;          �  ��       =             �       P          �   `                              ;          �  ��       =             ��       P          �   �                      �       �         �   y�       �             g�       (          �    f                       `       �              ~       �         �   �       (                �                             �          @   ��      @         �   �                 @    `                             �              ��      @         �   ��                      �                      �      `               y�      �         ,h    g�      
          �     f                       `      `         �    ~      �         ;�    �      
          @     �                            �         �    ��     �         ;�    �               @     �                      �     �         �          �         ;�                     @     ��                             �                �     �         ,h           �         �     ��      �                      �                �     �         �     �     �                ��      �                �      �               �      �         �     �     @               ��      @                �      H                �      �         �     �     @               ��      @                �               �    �      F         @           �         �    8��                                        �    ?                @    ?        �         �   ���                              2         �   ��                @   ��       l         �   8�                      8        1         �   ��       1         @   �       N         �   q�                       �         �        �   ��        �        @   ��                �  �                                  @        �  �?         �        @  ��                 �  p                        p                  �  ��        @           �8        q�        �  �                       �                  �  ���                    ���        n�        �                                   .�        � �~         *�          ��         U`        � 8�                        �          .�        � ?��          �          ?�p         _`        ��                                   .�        ���         *�        |��         U`        �8                        8           Q      |��          Q      ���          .�    ��|q�                     �           N�        ���          N�    ����          1�    ?� ���                                    4�       �~?            x   ?� � ��           �        �p                       p            s�|   |  �q�           ��|   |   �8            '���������                                      )����������            ?�������� ��             �|   |  �               �                       /���������~             ��������� �              ���������               ��������               ǃ��������p             ?�������� �               |   |  �                                       �        ��             ǃ��������               |   |   �                                        ?��������|               8|   |   �                        |                                        ���������               ���������               x                                                 ��   �                  ����                   �    �                                           �������                        �                  ������@                                           ~    �                        @                  ~    �                                                 �                                                 �                                                 `                                                 `                                   