�Ii  t�� �                                        <                     <                     <                     *                     r                     |                     ~                     *                     r                     |                     ~                     *                     r                     |                     ~                     *                     r                     |                     ~                     <                     <                                           <                     <                                          8                     <                     <                                          8                     <                     <                                          8                     <                  � <                                       � 8                     <                 ���<                                      ���8                     <               ������                                    ������                     <               �������                                    �������                     <              �������                                   �������                     <              ?�������                                   ?�������                     <             ��������                                  ��������                     <            ���������                                 ���������                     <            ���������                                 ���������                     <            ���������                                 ���������                     <            ����������                                 ����������                     <           ����������                                ����������                     <           ����������                                ����������                     <           ����������                                ����������                     <           ����������                                ����������                     <           ����������                                ����������                     <           ����������                                ����������                     <           ����������                                ����������                     <           ����������                                ����������                     <           ����������                                ����������                     <           ����������                                ����������                     <           ����������                                ����������                     <           ����������                                ����������                     <           ����������                                ����������                     <           ����������                                ����������                     <           ����������                                ����������                     <           ����������                                ����������                     <           ����������                                ����������                     <           ����������                                ����������                     <           ����������                                ����������                     <          �����������                               �����������                     <          �����������                               �����������                     <          �����������                               �����������                     <          ������������                               ������������                     <         ������������                              ������������                     <        �������������                             �������������                     <        �������������                             �������������                     <       ��������������                            ��������������                     <       ?��������������                            ?��������������                     <     ����������������                          ����������������                     <  �������������������                       �������������������                     <  ��������������������                       ��������������������                     <  �������������������                       �������������������                     <  ?�������������������                       ?�������������������                     <  �������������������                       �������������������                     <  �������������������                       �������������������                     <  �������������������                       �������������������                     <   �������������������                        �������������������                     <   ������������������                        ������������������                     <   ������������������                        ������������������                     <   ������������������                        ������������������                     <   ������������������                        ������������������                     <   ������������������                        ������������������                     <    �����������������                         �����������������                     <    �����������������                         �����������������                     <    �����������������                         �����������������                     <    �����������������                         �����������������                     <     ?�������  <������                         ?�������  <������                    <     �������   �����                         �������   �����                    <     �������    C����            |             �������    C����            |        <      ������     ?���            |              ������     ?���            |        <      ������     ���            |              ������     ���            |        <       ������      ��                           ������      ��                    <       �����      ��                           �����      ��                    <        {����       ��                            {����       ��                    <         ����       �                              ����       �                     <         ���       �                              ���       �                     <                    �                                         �                     <                     |                                          x                     <                     <                                          8                     <                     <                                          8                     <                     <                                          8                     <                     <                                          8                     <                     <                                          8                     <                     <                                          8                     <                     <                                          8                     <                     <                                          8                     <                     <                                          8                     <                     <                                          8                     <                     <                                          8                     <                     <                                          8                     <                     <                                          8                     <                     <                                          8                     <                     <                                          8                     <                     <                                          8                     <                     <                                          8                     <                     <                                          8                     <              ������<              ������              ������8              ������<                   <              ������              ������8              ������<              �����<              �                  ������8              ������<              �����<              �                  ������8              ������<              �����<              �                  ��DTG�8              ��DTG�<              �����<              �                  ���U��8              ���U��<              �����<              �                  ���U��8              ���U��<              �����<              �                  ���L��8              ���L��<              �����<              �                  ���U��8              ���U��<              �����<              �                  ���U��8              ���U��<              �����<              �                  ���TG�8              ���TG�<              �����<              �                  ������8              ������<              �����<              �                  ������8              ������<              �����<              �����              �   �8              ������<              �  �<              ��                �   �8              ��  �<              �  �<              ��                �   �8              ��  �<              �  �<              ��                �   �8              ��  �<              �  �<              ��                �   �8              ��  �<              �  �<              ��                �   �8              ��  �<              �  �<              ��                �   �8              ��  �<              �  �<              ��                �   �8              ��  �<              �  �<              ��                �   �8              ��  �<              �  �<              ��                �   �8              ��  �<              �  �<              ��                �   �8              ��  �<              �  �<              ��                �   �8              ��  �<              �  �<              ��                �   �8              ��  �<              �  �<              ��                �   �8              ��  �<              �  �<              ��                �   �8              ��  �<              �  �<              ��                �   �8              ��  �<              �  �<              ��                �   �8              ��  �<                 �<              �����              ������8              ������<              �����<              �                  ������8              ������<                   <                                 ������8              ������<              ������<              ������                     8              ������<                  � <                9 �                 > � 8                ? � <            �����������          �����������          �����������          �����������                               �����������          �����������          �����������          �����������                               �����������          �����������          �����������                               �����������          �����������          �����������                               �����������          �����������          �����������                               �����������          �����������          �����������                               �����������          �����������          �����������                               �����������          �����������          �����������          ?���������           �����������          �����������          �        �          ?���������           �����������          �����������          ����������          0                   �����������          �����������          �����������          7���������           �        7�          �        ?�          �����������          4        H           �        7�          �        ?�          �����������          4        H           �        7�          �        ?�          �����������          4        H           �        7�          �        ?�          �����������          4        H           �        7�          �        ?�          �����������          4        H           �        7�          �        ?�          �����������          4     0 H           �     0 7�          �     0 ?�          �����������          4     � H           �     � 7�          �     � ?�          �����������          4 ��`� H           � ��`� 7�          � ��`� ?�          �����������          4�����?�H           ������?�7�          ������?�?�          �����������          4����� H           ������ 7�          ������ ?�          �����������          4����� H           ������ 7�          ������ ?�          �����������          4����� H           ������ 7�          ������ ?�          �����������          4����� H           ������ 7�          ������ ?�          �����������          4����� H           ������ 7�          ������ ?�          �����������          4����� H           ������ 7�          ������ ?�          �����������          4����� H           ������ 7�          ������ ?�          �����������          4���� H           ����� 7�          ����� ?�          �����������          4� ��� H           �� ��� 7�          �� ��� ?�          �����������          4� ��� H           �� ��� 7�          �� ��� ?�          �����������          4� ��p H           �� ��p 7�          �� ��p ?�          �����������          4�      H           ��      7�          ��      ?�          �����������          4�      H           ��      7�          ��      ?�          �����������          4�      H           ��      7�          ��      ?�          �����������          4�      H           ��      7�          ��      ?�          �����������          4�      H           ��      7�          ��      ?�          �����������          4�      H           ��      7�          ��      ?�          �����������          4        H           �        7�          �        ?�          �����������          4        H           �        7�          �        ?�          �        /�          7���������           �        7�          �        ?�          ����������          0                   �����������          �����������          �        �                              �����������          �����������          �����������          ?���������           �        �          �����������          �����������                               �����������          �����������          �����������                               �����������          �����������          �����������          ?���������           �       �          �����������          �����������              �              ����������          �����������          �����������              �              ����������          �����������          �����������              �              ����|�����          ����������          �����������              �              �����|�����          �����������          �����������              �              �����x����          ����������          �����������              �              ��cxppL?�          ��c�ppL?�          �����������              �              �3&d�s1&I��          �3&d��1&I��          �����������              �              ��&|s3&H�          ��&|�3&H�          �����������              �              ��&|�p3&I��          ��&|��3&I��          �����������              �              ��&d�g�&I��          ��&d��&I��          �����������              �              ��gg�0L?�          ��g�0L?�          �����������              �              ���������          ����������          �����������              �              ����������          �����������          �����������              �              ����������          �����������          �����������              �              ����������          �����������          �����������              �              ����������          �����������          �����������              �              ����������          �����������          �����������              �              ����������          �����������          �����������              �              ����������          �����������          �����������              �              ����������          �����������          �����������              �              ����������          �����������          �����������              �              ����������          �����������          �����������              �              ����������          �����������          �����������           c`�x��           ����������          �����������          �����������           c �͛           ����������          �����������          �����������           c ��           ����������          �����������          �����������           cg���           ����������          �����������          �����������           l݂�9�           ����������          �����������          �����������           clق��           ����������          �����������          �����������           clق��           ����������          �����������          �����������           clق�͛           ����������          �����������          �����������           cgق�x��           ����������          �����������          �����������             ��              ����������          �����������          �����������            ��              ����������          �����������          �����������              �              ����������          �����������          �����������              �              ����������          �����������          �����������              �              ����������          �����������          �����������              �              ����������          �����������          �����������              �              ����������          �����������          �����������             � p            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������           ���S�           ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������           ���S�           ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������           ���S�           ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������           ���S�           ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������           ���S�           ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������           ���S�           ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������           ���S�           ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������           ���S�           ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������           ���S�           ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������           ���S�           ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � P            ����������          �����������          �����������             � p            ����������          �����������          �����������              �              ����������          �����������          �����������              �              ����������          �����������          �����������              �              ����������          �����������          �����������              �              ����������          �����������          �����������              �              ����������          �����������          �����������             � �            ����������          �����������          �����������             ��            ����������          �����������          �����������             ��            ����������          �����������          �����������           fb��            ����������          �����������          �����������           3fb��            ����������          �����������          �����������           3?�            ����������          �����������          �����������           3?�            ����������          �����������          �����������           3���            ����������          �����������          �����������           ��� �            ����������          �����������          �����������              �              ����������          �����������          �����������              �              ����������          �����������          �����������              �              ����������          �����������          �����������              �              ����������          �����������          �����������              �              ����������          �����������          �����������              �              ����������          �����������          �����������              �              ����������          �����������          �����������              �              ����������          �����������          �   �   �          ?���������           ����������          �����������          �����������                               �����������          �����������          �����������                               �����������          �����������          �����������                               �����������          �����������          �����������                               �����������          �����������          �����������                               �����������          �����������                                                    �����������          �����������          �����������          �����������                                �����������                   <                     <                                           <                     <                                          8                     <                     <                                          8                     <            �����������          �����������          �����������          �����������                               �����������          �����������          �����������          �����������                               �����������          �����������          �����������                               �����������          �����������          �����������                               �����������          �����������          �����������                               �����������          �����������          �����������                               �����������          �����������          �����������                               �����������          �����������          �����������                               �����������          �����������          �����������                               �?�?�������          �?�?�������          �����������                               �?�?�������          �?�?�������          �����������                               �?�������          �?�������          �����������                               � �13�0q��          � �13�0q��          �����������                               �"I32dɑ$��          �"I32dɑ$��          �����������                               �&g32|ɓ3��          �&g32|ɓ3��          �����������                               �&s32|ɓ9��          �&s32|ɓ9��          �����������                               �&I3"dɓ$��          �&I3"dɓ$��          �����������                               �&c��L31��          �&c��L31��          �����������                               �����������          �����������          �����������                               �����������          �����������          �����������                               �����������          �����������          �����������                               �����������          �����������          �����������                               �����������          �����������          �����������                               �����������          �����������          �����������                               �����������          �����������          �����������                               �����������          �����������                                                    �����������          �����������          �����������          �����������                                �����������                   <                                          8                     <                     <                                          8                     <                     <                                          8                     <            �����������          �����������          �����������          �����������                               �����������          �����������          �����������          �����������                               �����������          �����������          �����������                               �����������          �����������          �����������                               �����������          �����������          �����������                               �����������          �����������          �����������            ������             �����������          �����������          �����������            �                 �����������          �����������          �����������            �                 �����������          �����������          �����������            �                 �����������          �����������          �����������            �                 �����L����          �����L����          �����������            �                 ���ϞO?����          ���ϞO?����          �����������            �                 ������?����          ������?����          �����������            �                 ������?����          ������?����          �����������            �                 ������?����          ������?����          �����������            �                 ������?����          ������?����          �����������            �                 ������?����          ������?����          �����������            �                 ���ϞO?����          ���ϞO?����          �����������            �                 �����O?����          �����O?����          �����������            �                 �����������          �����������          �����������            �                 �����������          �����������          �����������            �                 �����������          �����������          �����������            ������             ��     ���          �����������          �����������                               �����������          �����������          �����������                               �����������          �����������          �����������                               �����������          �����������                                                    �����������          �����������          �����������          �����������                                �����������          �����������          �����������                                �����������