�;`  �82]         �0     �  �   ` 0                   �0     �  �   ` 0                   �0     �  �   ` 0                   �0     �  �   ` 0                   �0    �  � ` ` 0                   �0    �  � ` ` 0                   �0    �  � ` ` 0                   �0    �  � ` ` 0                    0    �  � ` ` 0                    0    �  � ` ` 0                    0    �  � ` ` 0                    0    �  � ` ` 0                   3ǜ>̓�|�sl�Ǐ3�                  3ǜ>̓�|�sl�Ǐ3�                  3ǜ>̓�|�sl�Ǐ3�                  3ǜ>̓�|�sl�Ǐ3�                  ��l��m�v�cm��ٶl                  ��l��m�v�cm��ٶl                  ��l��m�v�cm��ٶl                  ��l��m�v�cm��ٶl                   ߷��m�f�cm���l                   ߷��m�f�cm���l                   ߷��m�f�cm���l                   ߷��m�f�cm���l                                                                                                 �6�m�3f�cm���l                                                                                                                                       ٶl��m�3f�a͛ٶl                                                                                                                                       �3ǌ�́�f�1���3��                                                                                                                                                    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 �                           �        �              0            �        �                                     �             <            �       �    0         <            �       �    8         8            ��       �             8             �        �             :            �        |�   6         9            ��       |�   >         >            ��       ?��            8                    <�   �        ;�           �        ���   3�        8�           7��       ���   ?�        ?�           ?��       ��            8�                    s��   �        ;�           ��      ���   7�        8�           o��      ���   ?�        ?�           ��       ���            8�            @       ���   x        ;�           ?��      ��p   3�        8�           ���      ��p   ?�        ?�           ���      ���            8�                    ��p   �        ;�          ��      ���   7�        8�          ���      ���   ?�        ?�          ���      ���            8�           @        ���   �       ;�@          ���      ��   3��       8�@         ��      ��   ?��       ?��         ���      ���            8�           �        ��   ��       ;�         ��      ��   7��       8�         ���      ��   ?��       ?��         ���      ���            8�                    ��   �       ;�         ���      ���   3��       8�         ���      ���   ?��       ?��         ���      ���            8�                   ���   ��       ;�          ���      ���   7��       8�         ���      ���   ?��       ?��         ���      ���            8�                    ���   ��      ;� @        ���      ���   3���      8� @        ���      �F   ?���      ?���        ���      ���            8�                   �@   ���      ;�           ���      v,   7���      8�          ���      
���   ?���      ?���        ���      v<            8�           [              ��      ;�           �_�      ��   3���      8�          ���      �n�   ?���      ?���        �z�      �0            8�                           ���      ;�           ���      ���   7���      8�          ���      ���   ?���      ?���        ���                    8�                           ��      ;�           ���      ���   3���      8�          ���      ���   ?���      ?���        ���      �            8�                     �    ���      ;�          ��      wj�   7���      8�          ���      ��   ?���      ?���        ���       �j             8�                     j    ��      ;��@         ��      ��   3���      8ڠ@        ���      ��   ?���      ?���        ���       �     �       8��                          ��      ;��         ?��      ���   7��      8��@        ���      ���   ?��      ?��        ���       @ @            8�                           ��      ;�           ��      ��p   3���      8�           ���      ��p   ?���      ?���         ���         �            8�                           ��       ;� �         ��      ���   7��       8� �         ��      ���   ?��       ?��          ��                    8�                           �       ;�           ��       ���   3��       8� �         ?��       ���   ?��       ?��          ?��                    8�                           ��       ;�           �        |�   7��       8�           ��       |�   ?��       ?��          ��       �             8�                                                  ��       �                           ��       �                           ��                                                                                   �                           �        �                           �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          ��  �    0          �  �    ��                                                                                                                         �  ` �    1�          �  ��   ��                                                                                                                         �  ` �    00          �  ��   ��                                                                                                                         �y�s��    0>s���      ��|珀   ��                                                                                                                      ��fl�    0;fm�`      �v�ـ   ��3m�                                                                                                                      �}�g��    03fm��      ��f�ـ   ��3m�                                                                                                                      �ͳf�    03fm�       ��f��   ��3m�                                                                                                                      �ͳfl�    1�fm�`      ��f�ـ   ��3m�                                                                                                                      �}�3��    3cͳ�      ��fg��    ��m�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �                                    @                                                                                                                     �   c   �                �`� �   @                                                                                                                     �   c   �               � � �   @                                                                                                                     �   c   �               � � �   @                                                                                                                     �   c<�9���             ��o��<y�   @                                                                                                                     ����fͳm�6c����      �����nٳf�����                                                                                                                         cf�?1�7�              ��lٳ`}�                                                                                                                             cf�0�6               ��lٳ`̀                                                                                                                             cfͳm�6`              �slٳf̀                                                                                                                             c<�9���               �clϳ<}�                                                                                                                                                     `                                                                                                                                                          �                                                 