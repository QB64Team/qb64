��j  T��                        �    `�       �                                               �    `�       �                                               �    `�       �                                               �    `�       �                                               0   �� �     �                                               0   �� �     �                                               0   �� �     �                                               0   �� �     �                                                   �� �     �                                                   �� �     �                                                   �� �     �                                                   �� �     �                                               ����睰���<��<�8                                              ����睰���<��<�8                                              ����睰���<��<�8                                              ����睰���<��<�8                                              �m�6 `���6��0�3fٰ                                              �m�6 `���6��0�3fٰ                                              �m�6 `���6��0�3fٰ                                              �m�6 `���6��0�3fٰ                                                                                                                                                                                     7���������>͘0fٰ                                                                                                                                                                                                                                                        6�`����� f͘0fٰ                                                                                                                                                                                                                                                       6m�6`�ٰ6Û0f͘3fٰ                                                                                                                                                                                                                                                       �����Ǚ�c�>��<�3l                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �             �                                                  �             �                                                  �             �                                                  �             �                                                  �             �                                                  �             �                                                  �             �                                                  �             �                                                  �             �                                                  �             �                                                  �             �                                                  �             �                                                                                                                                                                                        �             �                                                                                                                     �             �                                                  �             �                                                  �             �                                                  �             �                                                                                                                 
                                                                                                                                                                                             <             <                                                
<             <                                                                                                                                                                          #             #                    �             �             #             #                    �             �             >             >                    �             �             "             "                    �             �             Lj             Nj                    `             `             Tj             Jj                    `             `             \6             \6                    �             �             H*             H*                    @             @             xF             tF                    @             @             xF             |F                    @             @             x|             p|                    �             �             pD             pD                    @             @             ��             ��                   �            �             ��             ��                   �            �             �|             �|                   �            �             �D             �D                   �            �             �             �                   ��            ��            ��            ��                   ��            ��             3�             3�                   ��            ��             3�             3�                   ��            ��             ��             ��                   �            �            ��            ��                   �            �             0�             0�                   �             �              0�             0�                   �             �              ��             ��                   �             �              ?�             ?�                   �             �              �0             �0                   �             �              00             00                   �             �             p�            p�                   �             �             ��            O�                   �             �             �<            �<                   �             �             @            @                   �             �              ��            ��                   ��            ��            C�            ��                   ��            ��            �2             �2                   ��            ��             �             �                   ��            ��            ��            ��                   ��            ��            H�            ��                   ~�            ~�            	�1            	�1                   ��            ��            �             �                     �             �            ��            O�                   f�            �            �            �                   ހ            ��            ��            �                   a�            a�                                             ��             �            �>            ��                   O             �             �            GL                   �             �             �2            ��                   I                                                           �                                      ��                   �                          .             ހ                   �             �             >                               �                                                                                       3             3��                   
�                           5.             2��                   �                           '>             '                    �                           "             "                    	                            (             ?                                  2              
\             �                    /                            |                                                                                               2                            f(             g                                  6              j\             e                    /              2              N|             N:                    =                            D              D                                                P             ~                    "              d              �             z                    ^              .              �             4                    :              0              @             0                    d                             �P             �>                    *              l              Ը             �:                    ^              d              ��             �t                    z              0              �@             �0                    $                             �             4�                    D              �              )p             >�                    �              \              9�             h                    t              `              �             `                    �              @             ��            �|                    T              �             �p            �t                    �              �             9�            8�                    �              `             �            `                    H              @              1@             i�                    �             �              R�             }�                   x              �              s�              �                    �              �              !               �                   �              �             1@            8�                    �             �             R�            (�                   x             �             s�            q�                   �              �             !              �                    �              �              b�             ��                                               ��             ��                   �             p              ��             A�                   �             �              B              A�                                               b�            q�                   P             `             ��            Q�                   �                           ��            �                   �             �             B             A�                                               �             ��                                 @             ˀ            ��                   �             �             π            �@                   �                           �             �                    @                           �             ��                   �             �             �            �                   �             @             o�            g@                   �                           d             c                    @                           �             ��                   @             �             �             �@                   �             �              ?              >�                   @                            8              >                    �                           �             ��                   '@             '�             �             �@                   ?�             ?�              ?              >�                   @                            >              >                    �                           ��            ��                   '�             '�             ��            ��                   ?�             ?�             =�            =�                   �             �              =�             =�                   �             �             ��             �                   �             �             �            ��                   ?�             ?�             �`             �                   �             �             <`             �                   �             �             |�            �                   �             7�             
�            ��                   /�             �             |0            |0                   �             1�             0            0                   !�             �             <�            �                   �             ?�             
G�            �                   +�             3�             |8            <8                   =�             �             $0            0                   �             �             V�            ~�                   #�             g�             ��            y�                   ^�             ,�             �0            60                   ;�             3�             @             0                    d�              �             Q�            ?�                   *h             l�             �`            
:`                   ^8             d8             ��            u�                   zh             0�             @             0                    $(              (             �`            4�`                   D              �              )p             >�                    �              \              9�`            h`                   t             `0             �             `                    �              @              �             |                    T              �              )p             t                    �              �              9�             8�                    �              `              �             `                    H              @              1@             i�                    �             �              R�             }�                   x              �              s�              �                    �              �              !               �                   �              �              1@             8�                    �             �              R�             (�                   x             �              s�             q�                   �              �              !               �                    �              �              b�             ��                                               ��             ��                   �             p              ��             A�                   �             �              B              A�                                                b�             q�                   P             `              ��             Q�                   �                            ��             �                   �             �              B              A�                                                �             ��                                 @             K�            ��                   �             �             π             �@                   �                            �              �                    @                            �              ��                   �             �             K�             ��                   �             @             π            �@                   �                            �              �                    @                           �             O�                   @             �             �             �@                   �             �             �             �                   @                                                            �                           �             ��                   @             �             �             G@                   �             �             �             ��                   @                                                            �                                        ��                   �                           .             ހ                   �             �             >                                 �                                                                                                     ��                   J�             K              .             ��                   ��             �              >                                 �                                                            	                            (             ?                    q              r              
\             �                    �              �              |                                                                                                B              @              (                                                             
\                                 �              �              |             :                                                                                                                 P             ~                                                �             z                    �              �              �             4                                                  @             0                                                  P             >                   @             @              �             
:                   ��            ��             �             t                    @              @              @             0                                                  �             4�                   �             �              )p             >�                   ߀            ߀             9�             h                                                  �             `                                                �             |                    0              0              )p             t                   �             �              9�             8�                                                  �             `                                                  1@             i�                                                R�             }�                   �             �              s�              �                                                  !               �                                                  1@             8�                                                R�             (�                   �             �              s�             q�                                                !               �                                                  b�             ��                   �             �              ��             ��                   ~             ~              ��             A�                    �              �              B              A�                                                b�             q�                    �              �              ��             Q�                   �             �              ��             �                                                  B              A�                                                  �             ��                    0              0             K�            ��                   �             �             π             �@                                                  �              �                                                   �              ��                                               K�             ��                   ;�             ;�             π            �@                                                �              �                                                  �             O�                                               �             �@                   -�             -�             �             �                                                                                                            �             ��                                               �             G@                   >�             >�             �             ��                                                                                                                             ��                    �              �             .             ހ                   ?p             ?p             >                                                                                                                                           ��                   P              P              .             ��                   ��             ��             >                                                                                                                            (             ?                    x              x              
\             �                    ��             ��             |                                                                                               @              @              (                                                             
\                                 ��             ��             |             :                                                                                                                  P             ~                                                �             z                    ��             ��             �             4                                                  @             0                                                  P             >                   @             @              �             
:                   ��            ��             �             t                    @              @              @             0                                                  �             4�                   �             �              )p             >�                   ߀            ߀             9�             h                                                  �             `                                                �             |                    0              0              )p             t                   �             �              9�             8�                                                  �             `                                                  1@             i�                                                R�             }�                   �             �              s�              �                                                  !               �                                                  1@             8�                                                 R�             (�                   �             �              s�             q�                                                !               �                                                  b�             ��                   �                            ��             ��                   ~             �              ��             A�                   �                            B              A�                                                b�             q�                   `                            ��             Q�                   �             |              ��             �                   �             �              B              A�                                                �             ��                   H             @             K�            ��                   �             �             π             �@                   �                            �              �                                                 �              ��                                 �             K�             ��                   �             `             π            �@                   �                            �              �                    @                           �             O�                   
�             �             �             �@                   �             �             �             �                   �                                                            @                           �             ��                                 �             �             G@                   �             �             �             ��                   @                                                            �                                        ��                                 	@             .             ހ                   �             �             >                                 @                                                            �                                        ��                                 �             .             ��                   3�             	�             >                                 �             <                                               -                            (             ?                    *              �             
\             �                    7�             �             |                                 >�             8                                                	                            (                                                             
\                                 g                            |             :                    =              x                                                Z                            P             ~                    T              %              �             z                    o              /              �             4                    }              p              @             0                                                 P             >                    0              .              �             
:                    �              &              �             t                    z              �              @             0                    �                             �             4�                    �              J              )p             >�                    �              ^              9�             h                    �              �              �             `                    $              @              �             |                    `              \              )p             t                   �              L              9�             8�                    �             �              �             `                   h              @              1@             i�                   P              �              R�             }�                   �              �              s�              �                   �             �              !               �                    H              �              1@             8�                    �              �              R�             (�                   8              �              s�             q�                   �             �              !               �                   �              �              b�             ��                   �             (              ��             ��                   x             x              ��             A�                   �             �              B              A�                    �                            b�             q�                   �             p              ��             Q�                   p             0              ��             �                   �             �              B              A�                   �                            �             ��                   @             P             K�            ��                   �             �             π             �@                   �                            �              �                                                 �              ��                                 �             K�             ��                   �             `             π            �@                   �                            �              �                    @                           �             O�                   
�             �             �             �@                   �             �             �             �                   �                                                            @                           �             ��                                 �             �             G@                   �             �             �             ��                   @                                                            �                                        ��                                 	@             .             ހ                   �             �             >                                 @                                                            �                                        ��                                 �             .             ��                   3�             	�             >                                 �             <                                               -                            (             ?                    *              �             
\             �                    7�             �             |                                 >�             8                                                	                            (                                                             
\                                 g                            |             :                    =              x                                                Z                            <P             :~                    T              %              <�             ?z                    o              /              �              4                    }              p               @              0                                                 |P             ~>                    0              .              |�             ~:                    �              &               �              t                    z              �               @              0                    �                             ��             ��                    �              J              �p             ��                    �              ^              9�             8h                    �              �              8�             8`                    $              @             8��            8��                    `              \             ;��            ;��                   �              L              80             8(                    �             �              8              8                    h              @             D�             D�8                   �                           ��            ��                   �              �              8              8                                               8              8                                                 �}�            �}�                   �              �             ���            ���                   �             �             8�            8�                    �             �             8�            8�                   �              �             �=�            �=�                   �              �             ���            ���                   �             �             8�            8�                   �             �             8�            8�                    �              �             ��            ��                   �              �             ���            ���                   �             �             8�            8�                   �             �             8�            8�                   �              �             D             D                    �                          ��            ��                   �             �                                                                                                                                              8�            8�                                 �             ;��            ;��                   �             `                                                  �                                                                 @                                                                 �              �                                                   �             �                                                   �                                                                                                                                                   �                                                                  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �          �             �0   � �   �0   � �                                                                                                                                                                                                              3     `      3     l              0      `    0      l                                                                                                                                                                                                              0     `      0                   0      `    0                                                                                                                                                                                                                    0|����g��     0|��������         3�<��>g��  3�<��>����                                                                                                                                                                                                          f��6l�۶     f��6lٛm�         �m�fͻf�۶  �m�fͻfٛm�                                                                                                                                                                                                          f͛7��6     f͛7�ٛm�         ��0fͳf�6  ��0fͳfٛm�                                                                                                                                                                                                          f͛6�6     f͛6ٛm�         60fͳf�6  60fͳfٛm�                                                                                                                                                                                                          3f͛6l�6     3f͛6llٛm�         �m�fͳf�6  �m�fͳflٛm�                                                                                                                                                                                                          |͙���3     |͙�����l�         3�<��>�3  3�<��>���l�                                                                                                                                                                                                           `  0           `  0                      �             �                                                                                                                                                                                                                  ` �           ` �                      � |            � |                                                                         