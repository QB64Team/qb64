��i  �}��                       �                                                     �                                                     �                                                     �                                                    3 � `   00                                               3 � `   00                                               3 � `   00                                               3 � `   00                                               0 � `   00                                               0 � `   00                                               0 � `   00                                               0 � `   00                                               0<�p<�8;s�s|�                                          0<�p<�8;s�s|�                                          0<�p<�8;s�s|�                                          0<�p<�8;s�s|�                                          fٳ`�ݰ3f`��                                          fٳ`�ݰ3f`��                                          fٳ`�ݰ3f`��                                          fٳ`�ݰ3f`��                                          ~߰`>�ٰ3g�c�                                          ~߰`>�ٰ3g�c�                                          ~߰`>�ٰ3g�c�                                          ~߰`>�ٰ3g�c�                                                                                                                                                              `�0`f�ٰ3f 31�                                                                                                                                                                                                                        3fٳ`f�ٰ3f`�a�                                                                                                                                                                                                                        <�0>Ǚ�c�s|�l                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��            ��            ��            ��                                                                                                                                                                                       �"|           �"|           �"|           �"|          ݀            ݀            ݀            ݀          "             "             "             "                                                                    /���          /���          /���          /���        � \           � \           � \           � \                                                                                                                             c�"~0          c�"~0          c�"~0          c�"~0        ݁�          ݁�          ݁�          ݁�        "           "           "           "                                                                  �/���         �/���         �/���         �/���        A� \          A� \          A� \          A� \                                                                                                                           s���s�        s���s�        s���s�        s���s�      �  �         �  �         �  �         �  �                                                                                                           3�����`        3�����`        3�����`        3�����`      `   1�        `   1�        `   1�        `   1�          @             @             @             @                                                                 �����        �����        �����        �����       �   @         �   @         �   @         �   @                                                                                                                 �������       �������       �������       �������      f    0        f    0        f    0        f    0                                                                                                                         o�����v       o�����v       o�����v       o�����v      �     �        �     �        �     �        �     �          D            D            D            D                                                               ��� ��       �������       �������       �������       �� &             &             &             &                                                                                                                         ��  ���      ��������      ��������      ��������    @ � x        @            @            @           �             �             �             �                                                                    >��   ���      >��������      >��������      >��������                                                           �             �             �             �                                                              m��   ?��      m��� ����      m��������      m��������        �@        �  @            @            @                                                                                                                        ���   �X      ���  ��X      ��������X      ��������X    ( `   0 �      (  � �  �      (       �      (       �                                                                                                               ��    ��     ���  ���     ���� ����     ���������    �    @           @        �   @             @    @             @             @             @                                                                    �     ��     ��   ?��     ��� ���     ��������    �           �   �       �  x �        �                                                                                                                              ��     �     ���   ��     ���  ���     ���������   @     �     @ `   0      @ �        @                                                                                                                              �     ?�     �    ��     ��   ��     ��� ����    �     @      � �          �   �       �  �                                                                                                                  ��     ��    ��    ���    ���   ���    ���� ����   `     0                  0   `         x �      �             �             �             �                                                                    �      �@    ��     ��@    ��    ��@    ���  ���@  	 �     �    	      �    	  �    �    	  �   �                                                                                                                      5�      �`    5��     �`    5��    ��`    5���   ��`  
      �    
      ��    
      �    
    � �           @             @             @             @                                                            /�      ��    /��     ?��    /��    ���    /���   ?���         @          @ @           @         @  @                                                                                                              [�       ��    [��     ��    [��     ��    [���   ���  $           $             $     �     $  `   0                                                                                                                        ��       �X    ���     �X    ���     ?�X    ���    ��X  (       �    ( @      �    (      @ �    (  �     �  @              @              @              @                                                                      ��       �    ��      ��    ���     ��    ���    ���  @       �@    @ �      @    @         @    @       @                                                                                                             o�       ?�   o�      ��   o��     ��   o��    ���  �       @     �            � @           �                    @              @              @              @                                                           _�       �   _�      ��   _��     ��   _��     ���  �              �            � @           �                                                                                                                             ��       �   ��       ��   ��      ��   ���     ��                              �                 �                                                                                                                  ��       �   ��       ��   ��      ��   ���     ?��  @                                       @   @              @              @              @                                                                     ��       �   ��       �   ��      ��   ���     �� @@           @       �    @           @                                                                                                                                       �   �       ?�   �      ��   ��     �� ��           �       @    �           � @                                                                                                                                    �   �       ?�   �       ��   ��     ��  ��           �       @    �           � @                                                                                                                       �        ��  ��       ��  ��       ���  ��      ���                                     �        �              �              �              �                                                                     
�        ��  
��       ��  
��       ��  
��      ���                                  �                                                                                                                                  
�        ��  
��       ��  
��       ��  
��      ���                                  �                                                                                                                                  �        ��  ��       ��  ��       ?��  ��      ���              @                   @                                                                                                                             �        ��  ��       ��  ��       ?��  ��      ���
            
 @           
        @    
                                                                                                                              �         ��  �        ��  ��       ?��  ��      ���
            
 �           
        @    
                                                                                                                              �         ��  �        ��  ��       ��  ��       ���
            
 �           
              
                                                                                                                              �         �@  �        �@  ��       �@  ��       ��@         �    �       �             �           �
              
              
              
                                                                      �         ��  �        ��  ��       ��  ��       ���
            
 �           
              
                                                                                                                              +�         �  +�        ��  +��       ��  +��       ���         �    �                                                                                                                                                       +�         �  +�        ��  +��       ��  +��       ��         �                @                   �                                                                                                                      ?�         ~�  ?�        ��  ?��       ��  ?��       ��          �@           @    @       @           �@                                                                                                                +�         �  +�        ��  +��       ��  +��       ��         �                @                   �                                                                                                                      +�         �  +�        ��  +��       ��  +��       ��         �                @                   �                                                                                                                      +�         �  +�        ��  +��       ��  +��       ��         �                @                   �                                                                                                                      ?�         ~�  ?�        ��  ?��       ��  ?��       ��          �@           @    @       @           �@                                                                                                                +�         �  +�        ��  +��       ��  +��       ��         �                @                   �                                                                                                                      +�         �  +�        ��  +��       ��  +��       ��         �                @                   �                                                                                                                      +�         �  +�        ��  +��       ��  +��       ��         �                @                   �                                                                                                                      ?�         ~�  ?�        ��  ?��       ��  ?��       ��          �@           @    @       @           �@                                                                                                                +�         �  +�        ��  +��       ��  +��       ��         �                @                   �                                                                                                                      +�         �  +�        ��  +��       ��  +��       ���         �    �                                                                                                                                                       �         ��  �        ��  ��       ��  ��       ���
            
 �           
              
                                                                                                                              �         �@  �        �@  ��       �@  ��       ��@         �    �       �             �           �
              
              
              
                                                                      �         ��  �        ��  ��       ��  ��       ���
            
 �           
              
                                                                                                                              �         ��  �        ��  ��       ?��  ��      ���
            
 �           
        @    
                                                                                                                              �        ��  ��       ��  ��       ?��  ��      ���
            
 @           
        @    
                                                                                                                              �        ��  ��       ��  ��       ?��  ��      ���              @                   @                                                                                                                             
�        ��  
��       ��  
��       ��  
��      ���                                  �                                                                                                                                  
�        ��  
��       ��  
��       ��  
��      ���                                  �                                                                                                                                  �        ��  ��       ��  ��       ���  ��      ���                                     �        �              �              �              �                                                                             �   �       ?�   �       ��   ��     ��  ��           �       @    �           � @                                                                                                                               �   �       ?�   �      ��   ��     �� ��           �       @    �           � @                                                                                                                            ��       �   ��       �   ��      ��   ���     �� @@           @       �    @           @                                                                                                                               ��       �   ��       ��   ��      ��   ���     ?��  @                                       @   @              @              @              @                                                                     ��       �   ��       ��   ��      ��   ���     ��                              �                 �                                                                                                                  _�       �   _�      ��   _��     ��   _��     ���  �              �            � @           �                                                                                                                             o�       ?�   o�      ��   o��     ��   o��    ���  �       @     �            � @           �                                                                                                                              ��       �    ��      ��    ���     ��    ���    ���  @       �@    @ �      @    @         @    @       @                                                                                                                      ��       ��    ���     ��    ���     ?��    ���    ���                @                 @        �                                                                                                                           �       ��    ��     ��    ��     ��    ���   ���                                    �         `   0                                                                                                                         ;�      ��    ;��     ?��    ;��    ���    ;���   ?���                   @                     @                                                                                                                        /�      �`    /��     �`    /��    ��`    /���   ��`         �          � �           �        �  �                                                                                                                      �      ��    ��     ���    ��    ���    ���  ����    �                           �             �                                                                                                                           �     ��    �    ���    ��   ���    ��� ����   �`     0      �           � 0   `       �  x �                                                                                                                         ��     ?�     ��    ��     ���   ��     ���� ����         @       �             �         �                                                                                                                          ��     �     ���   ��     ���  ���     ���������          �         `   0          �                                                                                                                                          ��     ��     ���   ?��     ���� ���     ���������                     �           x �                                                                                                                                         ��    ��     ���  ���     ���� ����     ���������    @�          @           @  �         @                                                                                                                               ���   ��      ���  ���      ���������      ���������     `   0         � �                                                                                                                                                    ��   ?��      ��� ����      ��������      ��������         �           �                                                                                                                                                          7��   ��`      7�������`      7�������`      7�������`         �             �             �             �                                                                                                                        �  ���      �������      �������      �������     � � x         �             �             �                                                                                                                              ��� ��       �������       �������       �������        ��                                                                                                                                                                        ������z       ������z       ������z       ������z          �            �            �            �                                                                                                                         �������       �������       �������       �������                                                                                                                                                                                    ^������        ^������        ^������        ^������      !    @        !    @        !    @        !    @                                                                                                                          ?������        ?������        ?������        ?������          @             @             @             @                                                                                                                           ������        ������        ������        ������                                                                                                                                                                    �����         �����         �����         �����                                                                                                                                                                                      }����          }����          }����          }����        "           "           "           "                                                                                                                             ����          ����          ����          ����                                                                                                                                                                                      ���           ���           ���           ���          "             "             "             "                                                                                                                               ��            ��            ��            ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ?                                                                                                                                                                                                    3                          0             3                                                                                                                                                                                                                   0             0                                                                                                                                                                                         ���          ���          >���          0���                                                                                                                                                                                      훰          훰          3훰          >훰                                                                                                                                                                                      ̓0          6̓0          ̓0          3̓0                                                                                                                                                                                      ̓0          ?̓0          ̓0          3̓0                                                                                                                                                                                      3͛0          ͛0          3͛0          3͛0                                                                                                                                                                                      ��0          ��0          ��0          ��0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              