��V  ��0]                                            �������������������������            �������������������������                                                  �������������������������                                                                                      �������������������������            ?�������������������������            @                                    @                                    ?�������������������������            �������������������������            �                                    �                                    �������������������������            �                                   �������������������������           �������������������������            �                                   �                                   ��������������������������          ��������������������������          �                                   �                        �          '�������������������������@          '�������������������������@          �                        �          �                        �          G�������������������������           G�������������������������           �                        �          x                        �          ��������������������������          ��������������������������          x                        �          �                         �          !�������������������������          !�������������������������          �                         �          =�                         x          B��������������������������          B                        ?�          =�  ����   ����   ����   x          {�                         <          ���������������������������          �                        �          {�$�F�m��I$m��nI$�F�m��I <          ��                                  ?��������������������������                                  �          ��  ����   ����   ����            �                                  ���������������������������        @                        ��        �  ����   ����   ����            �                          �         ���������������������������@         �                        �@        �I$�F�m��I$m��nI$�F�m��I$�        �                          �        A���������������������������         A                         �         �   ����   ����   ����   �        |                          �        ����������������������������        �                          �        |   ����   ����   ����   �        �                           �        !���������������������������        !                                  �I$�F�m��I$m��nI$�F�m��I$ �        =�                           x        B����������������������������        B                          ?�        =�   ����   ����   ����   �x        {�                           <        �����������������������������        �                          �        {�   ����   ����   ����   �<        ��                                  ?����������������������������                                  �        ��I$�F�m��I$m��nI$�F�m��I$`        �                                  ����������������������������       @                          �        �   ����   ����   ����   �        �                                   �����������������������������       �                          �        �|   ����   ����   ����   �        �                                   �����������������������������                                  �        �nI$�F�m��I$m��nI$�F�m��I$l        �                                   �����������������������������                                   �        ��   ����   ����   ����   �        �                                   �����������������������������                                   q        ��   ����   ����   ����   ��        �                                   �����������������������������                                   1        䑶�m�$�Im�ےI$���m�$�Im�ےN        �                                   �����������������������������                                           �����   ?���   ����   ?���         �                                   �����������������������������                                           �����   ?���   ����   ?���         �                                   �����������������������������                                           䑶�m�$�Im�ےI$���m�$�Im�ےN        �                                   �����������������������������                                           �����   ?���   ����   ?���         �                                   �����������������������������                                           �����   ?���   ����   ?���         �                                   �����������������������������                                           䑶�m�$�Im�ےI$���m�$�Im�ےN        �                                   �����������������������������                                           �����   ?���   ����   ?���         �                                   �����������������������������                                           �����   ?���   ����   ?���         �                                   �����������������������������                                           䑶�m�$�Im�ےI$���m�$�Im�ےN        �                                   �����������������������������          >                                �����   ?���   ����   ?���         �   >                    �          ����������������������������          ��                   �           �����   ?���   ����   ?���         �   �                  d          ����������������������������         �@                  �           䑶���$�Im�ےI$���m�$�I��ےN        �   �                  �          ���������������������������         �                   �           �����   ?���   ����   ?���         �   A�                  �          ���A�������������������������         �                              �����   ?���   ����   ?���         �    `                  �         ��� ����������������������                            ��          䑶� y$�Im�ےI$���m�$�I��ےN        �    `                  ��         ��� �����������������������                            �          ��� p   ?���   ����   ?���         �                      ��         ��� ?����������������������                            �          ��� 0   ?���   ����   ?���         �                      �         ��� ����������������������                            �          䑶� $�Im�ےI$���m�$�I�ےN        �                      �         ��� ������������������� ���                            �          ���    ?���   ����   >��         �                                ��� ?�����������������������                                        ��� 0   ?���   ����   >��         �                      �          ��� ?������������������������                                        䑶� 9$�Im�ےI$���m�$�I��ےN        �                       �          ��� �����������������������          @                  �           ��� p   ?���   ����   ?���         �   �                    p          ����������������������������          ��                   �           �����   ?���   ����   ?���         �   >                               �����������������������������          >                                䑶��$�Im�ےI$���m�$�Im�ےN        �                                   �����������������������������                                           �����   ?���   ����   ?���         �                                   �����������������������������                                           �����   ?���   ����   ?���         �                                   �����������������������������                                           䑶�m�$�Im�ےI$���m�$�Im�ےN        �                                   �����������������������������                                           �����   ?���   ����   ?���         �                                   �����������������������������                                           �����   ?���   ����   ?���         �                                   �����������������������������                                           �nI$�F�m��I$m��nI$�F�m��I$m�        �                                   �����������������������������                                           ��   ����   ����   ����   ��        �                                   �����������������������������                                           ��   ����   ����   ����   ��        �                                   �����������������������������                                           �nI$�F�m��I$m��nI$�F�m��I$m�        �                                   �����������������������������                                   !        ��   ����   ����   ����   ��        x                            <       ������������������������������       �                            C        {�   ����   ����   ����   ��        <                            z       ������������������������������       �                            �        =nI$�F�m��I$m��nI$�F�m��I$mz                                    �       �����������������������������	       �                           	        �   ����   ����   ����   ��                                   �       �����������������������������       ��                                  |   ����   ����   ����   ��        �                          �       ����������������������������!       �@                          !        �I$�F�m��I$m��nI$�F�m��I$k�        �                          �       �?���������������������������A       �                           A        �   ����   ����   ����   ��        �                          ~       �����������������������������       �                          �        �   ����   ����   ����   �~         �                          �       ����������������������������       �                          !         �I$�F�m��I$m��nI$�F�m��I$^�         x                          =�       �����������������������������       ��                          B         x   ����   ����   ����   ��         <                          {�       �����������������������������       ��                          �         <   ����   ����   ����   {�                                   ��       ����������������������������       ��                                  I$�F�m��I$m��nI$�F�m��I$��                                  ��       ����������������������������       ���                                    ����   ����   ����  ��         �                        ��       ���������������������������        ��@                                  �  ����   ����   ����  ��         �                        ��       ��?�������������������������@       ��                         @         �$�F�m��I$m��nI$�F�m��I'��         �                        �       ����������������������������       ��                        �         �  ����   ����   ����  �          �                        ��       ���������������������������        �����                  ���           �  ����   ����   ����  ��          ���                  �����       ���  �������������������          ���  @                               ����m��I$m��nI$�F�m�������          ?���                  �����       ���  ?�������������������          ���                                  ?�������   ����   ���������          ���                  �����       ���  �������������������          ���                                 �������   ����   ���������             �                    ��        ���������������������������         �����                  !���              ��m��I$m��nI$�F�m��  ��             x                  <  ��        ���������������������������         �����                  C���              {����   ����   ����  ��             <                  z  ��        ?���������������������������         ?�����                  ����              =����   ����   ���z  ��                               �  ��        �����������������������	���         �����                 	���              �m��I$m��nI$�F�m��  ��                              �  ��        ��������������������������          ������                ���               ���   ����   ����  ��             �                �  ��        ����������������������!��� @        �����@                !��� @             ����   ����   ����  ��             �                �  �         �����?�����������������A��� �        �����                 A��� �             ĒIm�ےI$���m�$�G�  �              �                ~  �         ��������������������������         �����                ����              �  ?���   ����  ~  �               �                �  �          �������������������������          �����                !���               �  ?���   ����  �  �               x                =�  �          �������������������������          �����                B���               x�Im�ےI$���m�$�=�  �               <                {�  �          ?�������������������������          ?�����                ����               <  ?���   ����  {�  �                               ��  �          ������������������������          �����               ���                 ?���   ����  ��  �                              ��  �          ������������������������           ������              ���                Im�ےI$���m�$���  �               �              ��  �          �������������������� ���@          �����@               ���@               � ?���   ���� ��  �               �              ��             �����?���������������@����          �����               @����               � ?���   ���� ��                  �              �             ������������������������           �����              ����                �Im�ےI$���m�$��                   �              ��              �������������������� ���            �����              ! ���                 � ?���   ���� ��                   x              =��              �������������������� ���            �����              B ���                 x ?���   ���� =��                   <              {��               ?�������������������� ���            ?�����              � ���                 <Im�ےI$���m�${��                                  ���                 ����������������� ���              ���              ���                  ?���   ���� ���                                  ���                  �����������������                   ���                                   ?���   ���� ���                                  ���                  ����������������                   ��                                  Im�ےI$���m�$���                         ��      ���                  ?��������  ������                   ?��                                   ?��������� ���                         ���     ���                  ��������  �����                   ��                                   ?���������� ���                        �����    ���                  �������    ?����                    ��                                   Im��������m�$���                        �����    ���                  �������    ���� @                  ��              @                     ?����������� ���                       ��  ���   ��                   ������ ��  ��� �                  ��     ��      �                     ?����  ����� ��                        �� ���   ��                   ������ � � ���                   ��     � �                         Im��� ���m�$��                        ?�` ��?�   ��                    �������� ����                    ��    �� �                         ?���` ��?��� ��                        ��� ���   ��                    ���� 8� ����                    �    8� �                         ?���� ����� ��                       �?� �� ��  ��                    ?������ � ��                    ?�   �� �                        Io�?� �� ��$��                       �?� ��?�  ��                    ������ ����                    �   �� ��                        ?��?� ��?�� ��                       ?�?������  ��                    ����?���?�8��                     �   ?�  ?�8                         ?��?� ���� ��                       � ?������  �                    ��� ��?����@                    �   ��  ��  @                     I� ?�   ���$�                      � �������  �                     ������ � ���                    �  ��  ��|  �                      ?�     ��� �                       � ������?� �                     �����   x ��                     �  ��  ��� �                        ?�      �?� �                       � ��������� �                      �����    p�                      �  �   ��� p                       ���      �����                       ��������� �                      q��#�   	���                      q  #��  ��� �                       ���       ���                       ?>�������� �                      1����   `��                      1  ���  ��� �                       ��>       ���                       ��?������� � �                      � �   ��                        ��  ����                       ���        ���                      ����������  �                      � � ����                        ?�  ����                      ���         ��                      ���������� ��                      � ���                        �� ��� ��                      ���    �   ��                      ������������p                      !�  �  ��?�                      ! ��  �� ?��                      ���         �p                      ������������8                      #�8      ?��                      # 8��  ��� ��                      ���         �8                      <������������8                      C�|0    @ ��                      C |��  ��� ��                      <���         �8                      :?����������=�                      E��@    @ ��                      E �?��  ��� ��                      :��         =�                      z~ ����������~�                      ����   @ ��                      ����  ��� ��                      z�           ~�                      v������������~                      ��    �p���                      �����  ��    ��                      v�          ~                      ��������������                     	�� � � @A�                     	���  �  �A�                      ��           ?�                      ��������������                     �@ ���  !��                    �?�� ~   �!��                     ��           �                     ��������������                     �  p   ��                    ����   ���                    ��           �                     ��?��������������                    $/� ��� x|@                    $/���~    �x|@                    ��           ���                    ���������������                    $'� ��` �|@                    $'���~� � ��|@                    ��     �    ��                    ����������������                    HC� 0��  �>                     HC ��~ � ��>                     ��            ��                    �~��������������                    P�� �@� @�                     P� � ?� � ?��                     �~            ��                    ^������������� ��                    �  G�����                    �  � 8 � ��                    ^�     ~�      ��                    ^������ ��������                    �  x��<A  �                    �   �  ������                    ^�     �     ��                    �������> ?�����xp                    B  �q����!  ��                    B   p '����������                    ��    > 8    xp                    �������>������8p                    !D p&?��8� �ǈ                    !D     ?��8;���ǈ                    ��   �>�     8p                    {����� >������<8                    "� `���0�?��                    "�    ���������                    {�   >��  � <8                    =w������>�����8                    B� �#���
 ���                    B�   `��������                    =w�   �>�p    8                    :�������>�����^                    E ����  ��                    E   ���������                    :��   3�>�    ^                    z�������������                    �  	<��� � �                    �  �<�������                    z��   ���   �                    u�������;�����                    �?� |��?��@ �                    �?� �|��?� ?���                    u�   ���;   �                    �������=�����                   
?� ���?�`  4�                   
?� ����?� ���                    ��   ��=�  �                    ����� � �~�����                   � ���?��� Bx�                  p ����?����x�                   �    � �~`  ��                   ����� �?� �?�����                   � $������x�                  x 
������� x�                  �   �?� �0� ��                   ׁ���� s��������À                  (�"H��  �<@                  (~� ���  �� <@                  ׀   7 s����   �À                  �����O�������À                  (� `@P�?��<@                  (���?��?��� <@                  �    /�O���   �À                  ������>?���������                  P� ��?���0 �                   P��� ?����                    �    _�>?���   }��                  ����������������                  Q� �   ��� �                   Q���~   ��                     �    ������   ~��                  n�������� ������                  �� x0���  G                   �����x0���                      n   �����    8��                  ^��������=������                  �� ��A�?  _                   ����|�A�?�                     ^   �����=    ��                  ]�����y��=�~����q�                  � e��  ��X� �                   �����  ��  ?�                   ]�  �y��=�~�   q�                  ]���� �����q�����q�                  � �#  1� � ?�                   ����#  1�  �                   ]�   �����q��   q�                  ]���� ;���������q�                  ���   D�@ ?�                   �����   D�� �                   ]�   ;������@   q�                  ;���� w?��������9�                  �����"�@p?�                   �������"�� �                   ;�  w?�����`   9�                  ;�����n������?���9�                  �� ��  �                   ���� ��� �                   ;�  �n������    9�                  ;���������n�?���9�                  � 	$? � �?�  �                   ���? � �?�� �                   ;�  ������n�0   9�                  ;���������� ���9�                  � �$  � H�� �                   ���$ � H��@ �                   ;� �������    9�                  w���������� ����                  � (D  � D�� �                   ���D � D��� �                   w�  �������    �                  w�����w���݀����                  �  P�  � "� �                   ���� � "�� �                   w�  /�w����݀   �                  s�����o����/����                  �  ^�  � � �                   ���� � �� �                   s�  !�o�����(   �                  p?���6������������                  ��  _��� > �"                   ������� >� "                   p    6��������  ��                  p?���������������                  �� �� �� 	0
"                   ���?� �� 	0	� �"                   p   @��������  ��                  p?������{���������                  ��~ ��  @� 	
�"                   ���?�  C� 		��"                   p   @��������  ��                  `?������w��o������                  ����@  � �
�                    ��  ?�@ #� �	��                   `   @������o�  ��                  `������o��o������                  �� /��@ � �;                    �� ?�@ � �8��                   `   @������o�  ��                  `���������h�����                  �� A�@ � ��                    �� >�@ � ����                   `   �������h  ��                  `���������������                  �� AA�@`�O�                    �� >A�@`�O���                   `   ��������  ��                  `����0 `�������                  �� A@$�����O�                    �� >@$�����O���                   `   ��������  ��                  `�����?��������                  �� A@$���O�                    �� >@$�����O���                   `   ��������  ��                  `����  �������                  �� A@$���O�                    �� >@$�����O���                   `   ��������  ��                  `������?��������                  ��@I@$�`�O�$                   �� 6@$�`�O���                   `   ��������  ��                  `������������                  ���]� � O�t�                   ��@*� � O�#���                   ` @�������  �                  o������/��������                  �@@I� � H$�                   �  6� � H���                   o�  ��������   �                  o������7��������                  �@ A� $� H �                   �  >� +� H���                   o�  ��������   �                  o������;��������                  �@ A� D� H �                   �  >� K� H���                   o�  ��������   �                  o������?��������                  �@ A��� H �                   �  >��� H���                   o�  ��������   �                  o���������������                  �@ A�@�� H �                   �  >�@�� H���                   o�  ���������   �                  o���������`;����                  �@ A~@  � �� �                   �  >~@ � �����                   o�  �������`:   �                  o���������`����                  �@ /�@  � �� �                   �   @ � �����                   o�  _������`   �                  o���������`����                  � �@  � ��� �                   �    @ � �����                   o�  _������`   �                  w����������������                  � ~ �  � 	���                   � �   � 	����                   w�  _��������   �                  w����������������                  �/� �9  � 	?��                   � � 9  � 	?�� ��                   w�  _��������   �                  t?�������������                  ��  Q� � /� ��                   ����� � /�� �                   t   .�������   �                  p?���o��������                  �� _�� � A� �                   ������ � A�� �                   p    o�����  �                  p?���w����ݿ������                  �� _��    "@4 "                   ������    "@3�  "                   p    w����ݿ�  ��                  p���������������                  �� /�D    D�) "                   �����D    D�&�  "                   p   �������  ��                  x���������?������                  �� ��$    H�+� B                   �����$    H�%@  B                   x  ������?�  ��                  x��������n������                  �� 	'�    ��I  B                   �����    ��F�  B                   x   �����n�  ��                  ����?n�����������                  G���   �P  D                   G�����   �O�  D                   �   ?n������  ��                  ����w?���������                  G����  #��@p D`                  G������  #���  D`                  �  w?����`  ��                  �����;����� ���w�                  #�
 �   G��@  �`                  #��� �   G���  �`                  �   �;����� @  w�                  ���������t ����w@                  #� �  1�� �  ��                  #����  1��   ��                  �   �����t �  w@                  �����y��=� ����o@                  � e��  ��X� `��                  �����  ��   ��                  �   �y��=� �  o@                   ����x���߁������                  � ���A� ~�  y                   ���|��A� ~  9                    �  x���߁   ��                   ����������������                  	 _�0��<�  !                   	���_�0��<   ?!                    ��  �����    ��                   v���������������                  � �?�  ��� �"                   ���~?�  ��  "                    v�   �����    ��                   {����>?���������                  �� ������
0 �B                   ����?����� ~B                    {|   @>?���   ��                   ;����?��������                  ā `@_��?���D                   Ā��?���?��� �D                    ;~    ?���   ��                   =������������{�                  �A�"O��  a�$���                   �@� ���  a� � ��                    =�   0����   {�                   �����~ ?�> ����w�                  �@� '�����I����                   �@x 
ǁ����@����                    �  ~ ?�> ��  w�                   �������  �����                  �@� �?����� C�                   �@p ��?�������                    �   ��  `   ��                   �����|���������                  � p ��?�~`  7�                   �   ���?�~ ���                    ߀  |����   ��                   _�������������                  �� G�?�|�@ �                   � �G�?�| ?���                    _   ����    ��                   n?�������������                  ��� 	7�?�9 � �                    ��� �7�?�8����                     n    ����   ��               8   ��������������     p            �O� ���f  �                 8  �O�  ���a�����       p             �    0���   ��               |   �������o�������     �            �O� �+��
 �d@                |  �O�  `�����d@      �             �    ��`   ���               �   ���������������    �      �   �'� `��0� H@              �  �'�   ������H@     �      �    �   ���  ����             �   �����ǀ��������    �      � (� �'� pF8�� �@H�    Q         �  �'�    8�;���H�     �      � 8�  �    ǀ�    ?��   q     �  �   ������ �?�����o�   �      �� ��  �����!  @��   #     �  �  ��  p@'���������    �      ��  �    @ �8   ?o�  #     �  �    ������ ��������� ?� �      �� �� @x��<A  � @       �  �  ��  �  ������ @ ?� �      ��   �      �    ~���       ?�  ~    ����������������� �  �      �� �	�  G����! @       ?�  ~  �	� � 8 � �! @ �  �      ��   �      ~�     ����       � 8    w ���������������  �� p      �C� ���� �@� @" �  �     � 8  ��� � ?� � ?�" � �� p      �C�   w            ���   �     �      {����������������  ��8       ��� ��~� 0��  B �      ~�    ��~ ��~ � �B � ��8       ���   {�            ���  
     �  �  ;�������������w��  ��  �   ��	� ��<@ ��` �D     x�  ���< ��~� � ��D  ��  �   ��	�   ;À    �     w��     ��x���  =�������������{� ������    �
�  ��8  ��� �   4    ��x��� ��8 ��~    �� ������   ���   =��           {�  ���4    �y���  �������������w�  �����    �
?�  ��  p   ��   �@   �y��� �� ���   ���  �����    ����   ��           w�   ����@   ?�`
��  ���������������  ���?�   @�?� �@ ��� ?�  �/�    ?�`�� � ?�� ~   ��  ���?�   @���  ��           ��  �?���    �  �  �������������>��  ?� 8 ?�   ��?�@ �� � � � ��:Ā   �   | � ��  �  ��  ?�   >�   �?�?��  ��           >�� ��ŀ   �  �  �������������~��     ?�  ��	�  ?�    �p�� ��?�@   �   < ?� ���  ��   �      >x  ����  ��          ~�� ��?��    p  �  ������������ ���   �  ?�  	����?��   @ � �"?��   p  < ?���  ���  �   �  >x  	����� ��          ��� �"?���   � ��  |�������������  � ��  ����  ��    @ ~ �&�@@   �  � � ����  ���  ~  �  ?�  ���"   |         ���� �&D@@    � ��  ?�?�������������   � ��  ��&r�  ��G�    @ < �L�?�      �  � � G���  ���  <   �  �  ��r   �         ���� ��8       � ��  ��������������   � �� ��g*?�  ��/�       8���T�      �  G� � /���  ���  8   �  �� ��g*<@   �         �������Tx�      p ��  ��������������    � �� ��7�$o�  ���  �  � ��oH��      p  �� � ���  ��       � �� ��7�&l�  �         ?������oL��0  8 � �  �������������� p   �8  �?�gO�� ��� � `?  ��Ο��  8     @ � ��� ���  `  p     �8  �<~gNF�  O�     �  ����� �x�Μ��  | �   <  � ����������� � �   x  ��G�� ���� � �@ �?���  |      < � �?�  ��  �@ �      x  �>G��  �        ��� �0|��  | �     � ��������� � � �     ��F�3� ����    �@ �?��g   l      � ���  ��� @ �       �F�3�  � @       �� � '�"<�g  �8�  ǀ  � ��������y� � �p�  �  ������  ��@�   ��� �����   � �  ǀ�  ��  ���� ��    �  ��ҟ���� I� �       y�$� ��?��  �|�  �  ���������w� � ���  �  ���t��  ���>   	���� ����?�   �    ��  > �  ���� ��    �  ���t���  ��       w� � ��>�?� �|�  �   �������� � � ���  �  ����	O���� �   ���  ��������    � �      �����  �     � ��?�	O�  ?��       � � �'�����  |�  ��  �������� ?� �   �   � ������ ` ��� <   ��� ���� �       p� �      �����         � ������� I���      ?�$� �C�����8    ��  �������� �� �  p    �� �����L  ��� ?� �� ?�  ����2� �     �� �   <  ���         ��������L�  ?���    x �� � ����2��     �p  �?�?�����  �      �� �����  q�� ���� ��  �����8>       �p q   �� � �         �������p  ?�?�   ��� � �����8>�     �p   �ǀ����  �     > �� �����?� q�� 8�������  �����<       �p q   8� ��         �������?� ���ǀ  ��F�� �����<�      8   ?��� �?�  �    >   p �������� 1��������� �����ÿ��      8 1   ����         p����d���� ��?��� �?��� �����˿��     8   � � ���  �    >>  p ���`��  1������� �� ����?���       8 1   ����       >   p�{�` ��8 ��� � ����� �������p  �?�     ��� ���  � 8 �  8 �_D�?�  ��� ?���8 ?��  �澈    �?�       ?���8    8 @   8�D�?� ����� ���F�� 8�f>� 8 �?� p   ��� ?�   � 8 �  �8 ��J�   ��� ���� ���  �����     ?�       ����    8      8�J�  ����� ?� �� 8d��� 8 �?� �     ��� ��   � 8 � � 8 ��D���  ���� ~�� ���  ������  ?�         ~��     8     8�D�� �� ��� �� �� 8�����8<� �     ��  ���   � x�> � < ��`���  ���� ��  ���  ������� < @          ��      x �>  @ <<�G`�#� ��O��  ���F�� x�����G�<  � �     �������   �   � � ��p?���� ����      ��� ���~����    �  p                  @  � ���p?�s�� �� ������� �� ��������8 �  �      �����    � p �  � ���r�a��� �����    ��������������8 H                    p �   @ ��Gr��#�� ��  �����  ���������G��8 �   �      �����    � p �  � �?��3����� �����    ?���� ��g�����8                       p        �?�3���� ��I'�����$�F��p�g����8  �  p       ���     � p �  �  =�_#��� ������  ����� {d�G��� 8  �                    p @     8=�#��� ��   ����   ��p{�>G�� x    ��       ��      � �      @!�"p�	 ������  ������ �C��D��=�8     ��                p      x!�"qp� ��   ����   �� �C��D��=�x   ��                � �   �� @�� � �������������� ���<@7�8   ��                p   �� x�� � ��I$m��nI$�F�� ���4@7�x    ��                � �   � @���@�� �������������� ���΀'�8    ��                p   � x���@�� ��   ����   �� ���΀'�x p  �                � � �  �� @���� a �������������� �7��� �8    �                p    �� x���� o ��   ����   �� �7��@��  �  �� �              �� � �� �;����� !����������������w���~  C8     ��                p    �� �;���� /���I$m��nI$�F���w��~  _� �  �� �              �� � �� ?�_���� �������������������_�~  <     ��                x    �� <�_�S������   ����   �������� ?� � �� �              �� �8�� ;�����@`����������������'���� ��     ��                8  @ �� <��#��@`���   ����   ���'�G��.��?� ��> �� �              ����|�� ;����  0����������������?_��  ` �   ��                8�  �� <�S�� 0���I$m��nI$�F���<��� `?���>�� �              ����|�� ;���������������������������  ��                8� �� <��������   ����   ������?��p>� 9�              ����|�� s�G�7O�������������������n� �  � >               � ( �� |�G�H�?���   ����   ����:� �� ?� 9�              ��� 8� s��� ����������������0�> 8�  ?� >               �  � |���	 ?���I$m��nI$�F���0� 8� �   � q�              ���   ?� ���� ����������������"��@< �   � ~               �   ?� ���� ���   ����   ���"��@<��     � q�              ��       ����0������������������`�     � ~                      ����0���   ����   �����`����       �              ��       ������ �������������������� �       �                      ������� ����I$m��nI$�F����������       �              ��       ������ �������������������� �       �                      ������� ����   ����   ����������     À              ���     ���r� ������������������?� �      �               �      ����r�����   ����   ������7����      ��              ���      ��?
� ����������������~?�  �      �               �      ����?
�����I$m��nI$�F����~?���  �   �               � �� �   ��  �������������� ���  �  �   �               � �   ����� ��   ����   �� ������ �                  � �� �   � H�  �������������� �  ��  x �   �                � �   �� J�� ��   ����   �� �� ���� �   <               � �� �   x� M�  �������������� �� ��   �   ?�                < �   �� M�?� Im�ےI$���m�$� �� ���� �   |               � �� �   �� BM�   �������������� �� ���    �   �                > �   ��� BM� �  ?���   ���� � �� ��� ��?���   �               � � �  �?�  �   �������������� �     ��   ��                 �  ��?�� � ��  ?���   ���� � �  ��?���  �               � ���  �?�     �������������� �  
   ��  ��                ��  ��?�� �� Im�ےI$���m�$� �� 
��?�� �  �               � ���  �?�  B   �������������� �  �   � �  ��                ��  ��?�� B��  ?���   ���� � �� ����|                    � ?��    > 8�  �   �������������� ?�  	  8 �    ��                �    ?���� ���  ?���   ���� � ?�� 	?���>    > <               � ?�|    | x�     < �������������� ?�     x �    ?��                �    ����  ?�� Im�ےI$���m�$� ?��  ����   � <               � ?�?   � x�      < �������������� ?�      x ��   ���                �   ������  ���  ?���   ���� � ?��  �����  � x               � ��  ?� ��       x �������������� �       �  ��  ���                ��  ?�� ���  ���  ?���   ���� � ���  ?������  ��x               � ���  ?�����    �x �������������� ��    ��  ?�  �?�                 �  ?� ���  ��� Im�ےI$���m�$� ���  ?������� �     ?�����    � ��������     � �����    ���� ��    �  �����      �����      ����� ��������  ?����������� � �������������> �       �      � �|?���|���    > � ����� � ���� �|    |�  A������      ����      ������� ���������  ?����������� � ����������ǃ�����       0`      � ��������ǀ   �� ����� 0` ���� ��   ��  8����      �ϟ��      p����� ��������� Im��������m�$� ������������  ��       @      � ���  ?�����  �� ����� @ ���� ���  ?��  ���?�      �����      <���� ���������  ?����������� � ������������� �       �      � ����� ����� � ����� � ���� ����� �  �?� ��      ����       ��� ���������  ?����������� � �������������� �       �      � ����� ������ � ����� � ���� ����� �  �  ��      ����      �  ?�� ��������� Im��������m�$� ��������� �� ?�  �            � �� �  ?  �� ?�  � ����� ���� �� �  ?   �����      �����      �����  ���������  ?����������� � ��������  �     ?       �      �  ��     ~  �     ?  ������ ����  ��     ~   ������      ��{��      ������  �������   ?����������� �  ��������  ?��    �       �      �  �    �  ?��    �  ������ ����  �    �    ����       ��{��       �����   ?�������  Im��������m�$�  �������  ?��   �       	�      �  ��   �  ?��   �  ����� � ����  ��   �    ?����       ��{��       ����   ?�������   ?����������� �  �������  ��   �             �  ?��   �  ��   �  �����  ����  ?��   �    ����       �����       ����   �������   ?����������� �  ?�������  ��   �        �      �  ��   �  ��   �  �����   ����  ��   �    ����       �����       ����   �������  Im��������m�$�  �������  ��   �               �  ��   ��  ��   �  ����� � ����  ��   ��     ����       �����       ���    �������   ?����������� �  �������  ��� ��               �  ��� ��  ��� ��  ����� @ ����  ��� ��     ��        �����        ?��    �������   ?����������� �  �������   ��� ?��         `      �  ��� �    ��� ?��  ����� 0  ����  ��� �      ��        �����        ��     �������  Im��������m�$�  ������    �����         �      �   ������    �����   �����   ����   ������                 �����                �����    ?����������� �   ������    �����                 �   ?�����    �����   �����    ����   ?�����                 �����                �����    ?����������� �   ?�����    �����                 �   �����    �����   �����    ?����   �����                                       �����   Im��    6�m�$�   �����    �����                 �   �����    �����   ��������������   �����                                       �����    ?���   ���� �   �����     �����                 �   ����      �����   ��������������   ����                                         �����    ?���   ���� �   ����      ���                  �    ?���      ���    ��������������    ?���                                         ���    ��I$m��nI$�F��    ?���      ���                  �    ���      ���    ��������������    ���                                         ���    ��   ����   ��    ���       ?�                   �     �        ?�     ��������������     �                                           ?�     ��   ����   ��     �                             �                      ��������������                                                         ��I$m��nI$�F��                                    �                      ��������������                                                         ��   ����   ��                                    �                      ��������������                                                         ��   ����   ��                                    �                      ��������������                                                         ��I$m��nI$�F��                                    �                      ��������������                                                         ��   ����   ��                                    �                      ��������������                      ��������������                                    �                      ���������������                                                                                              ���������������                      ���������������                      @                                  @                                  ���������������                      ���������������                      @                                  @                                  ���������������                                                            ���������������                      ���������������                                                                                                  ���������������                      ���������������                                                                                                  ���������������                      ���������������                                                                                                  ���������������                      ���������������                                                                                                  ���������������                      ���������������                                                                                                  ���������������                      ���������������                                                                                                  ���������������                      ���������������                                                                                                  ���������������                      ���������������                                                                                                  ���������������                      ���������������                                                                                                  ���������������                      ���������������                                                                                                  ���������������                      ���������������                                                                                                  ���������������                      ���������������                                                                                                  ���������������                      ���������������                                                               ���������                         ���        ���                      ���        ���                         ���������                            ���������                         ���        ���                      ���        ���                         ���������                            ���������                         ���        ���                      ���        ���                         ���������                            ���������                         ���        ���                      ���        ���                         ���������                            ���������                         ���        ���                      ���        ���                         ���������                            ���������                         ���        ���                      ���        ���                         ���������                            ���������                         ���        ���                      ���        ���                         ���������                            ���������                         ���        ���                      ���        ���                         ���������                            ���������                                    @                                    @                            ���������                            ���������                                    @                                    @                            ���������                            ���������                                    @                                    @                            ���������                            ���������                                    @                                    @                            ���������                            ���������                                    @                                    @                            ���������                            ���������                                    @                                    @                            ���������                            ���������                                    @                                    @                            ���������                            ���������                                    @                                    @                            ���������                            ���������                                    @                                    @                            ���������                            ���������                                    @                                    @                            ���������                            ���������                                    @                                    @                            ���������                                                                  ���������                            ���������                                                                                                        ���������                            ���������                                                                                                        ���������                            ���������                                                                                                        ���������                            ���������                                                                                                        ���������                            ���������                                                                                                        ���������                            ���������                                                                                                        ���������                            ���������                                                                                                        ���������                            ���������                                                                                                        ���������                            ���������                                                                                                                                                                                                        