�
t  0C  ���>��00��>  ��@@��  ����  ���  �    ���   �� � ���G��6��?������?�������>��  �����        ���>��00��>"�"����EDED����ğ��"�2������  @��   �� � ���G��6��?������?�������>��  �����        ���>��00��>  ��AED���FG�Gď������������PP���
��#����h.�<���2r���8<|x���>�?�������>��  �����        ���>��00����  ����@@����@@�������������������� ����� ����@ ���� @����  ���� 0 ����� ����          ��������0�����0����p��28�>O�>o���W������������ꢿ��ǀǂ���P@�f��d �_�`0 ��/�� �>0�>�����          ��������0�����0����p��8�>p�> ��� �����ǂ�������������B���_��UP�V_�@#���?�� �>��>����o�          ��������0�����0����p��8�>p�> ��� �������� ���� ���A �G��G���O�@+���?�������>����o�          ��������0�����0����p��8�>p�> ��� �������� ���� ���@ �@�@ �@@  � � �>0�>����o�              } }   ������� ���������p�� �   �  �p    ��� ����� � ������ ������~���� �  �� ��   �7� �   ��rI� � ?������ �����ǀ ��� �  �� ���    � 8    ���� � ?������ ������   ���� �  �� ���   �      ��� �������������7��    �?� �  7�  ��� �  m��      �͵� ?�������������G�    ��(�  G�� ���� (���       ���� ~|���������c����    ���0b ��� ���� 0��|       >��������������#��     3�� " �� ����  m��       ������������� ��#��  �� "  � ����  ���         ������������� ?�#� � ���" ���������       ?��<�������������C�   @��B  �� ��� �=o��         ��8�����������/�pG�p    @ �?�F p�� ��� ?��9���         /�px?����������7�p���`    � ?��� ��� ��  ��y��         7�pt~����������{�8����    � ������ ��  ��u~          {�8��������������8�    �@�
���� ��  ���           ��8��������������� 8   ������ �� @ ���        @ ���������������|�  �� @�������  �   ����           |��������������"�� �  @C�"��� � >  �C���           ?���?������������$?�@ � :   !�$?�?���   �!���           �������������� H_�    ��H_�����    �����            �������������� HO� ��  	��HO ���|  �����          oy���������������  a0 @�x�� ���� � ?��xox            �^��������������� ���� ��8� �   � ��8^�            ����������������B  �� �B  � p � �����     ��     ������� ������B @���x� �B  � ��������     �    �{������| ������� �σ��B  ��   �@O������{�   @0| p    �w������|������p� �L��q�4 ���     ��pw����w�   �|�     p������@|������x �1���`��   ���������  @|�   x�������|������8  F?��? ?�   �?��?�������   9�|��    8�������|�?����  �?��?�"  ?@  �?��?�����@��   g�|�0    ��������<������>@ x��?�A   >  �x��?���� ��  ��<�   ؀�����<�w������ ������   ����� ���   �<�v   ������<�{������ �����@ h  ����� ?���   �<�{   ������ �������� $'���!  ��� ���� �     � ���  ������������� .I������� ������    6���a  ����� ����?����� D��  ���� ;�  ���     n ����0  ����� ��������� ����`�<� ��  �`�<��      _ ����  ������|�������� !@���` ����@����      ��|���   ���������=������ @> ��� ����@> ��      �����=�   �������@7����� �`?�1��  ������`?�1��      ���@6   p����|?���{����� ����
  ���������  8   �|?���z   @��������{������8 ��! �?�  �7��3�! �?  x�  ����{��    ��������������� 3�F0  cA  x���F0  c>  8�  ��������   ���� w����w�������@  �@�@x����@  �?  8�   w����w��   ���� ���������8'�� D ��x���� D @8�  ������ @ ���� ���������� (�" �$�@@8���" �$�� �   �������@   ����������݀���  H~$ �"�@ 8��~$ �"�� �  7������݀`   ���������n ?���  PH   ���@ 8��H   ��ʀ � /�����n "   �����w����v ?���  "P�   ���  8���   ���� �  /�w����v     ����������� ���@  �	   D��  ?�� 	   D��� �  _�������    ����������� _���@  �	    $��  ?��<	    $��� �  C������� P   ���m�����݃����� @��  "|(����?�  "|'�    @m�����݃�   �������������� A�@ `>����@ `��   ��������  �����z����������A�@ �  ����@ �  �?�   ���������  ���������������� A 	 � �  � G 	 ��   ��������  ���������ߏ���� _� !  	 v    � '  	 p��   ������߈   ��� ��������� ��� @ 	/�   |�� @ 	/���   ������   ���|7�����`���� ��Ȁ����   |�Ȁ������  |7�����`   �����` ��`���� ��I������   |�I��������  �������`   �����?���`���� ��I����   |�I��������  �������`   �����  @�`���� ��I����   |�I��������  �������`   �����?���`�������I ����H  l�I ������  �������`   ��� 6���?��`��������  @ ��� �T��  � ��G�� � 6������`@ ��� 6���_��o���������  )  �
H  l��  '� ���   6������o�   ��� 6���o��o����� ���  I� �
   |��  W� ���   6������o�   ��� 6��zw��o����� ���  �� �
   |��  �� ���   6������o�   ��� 6�����o����� ��� 	� �
   |�� � ���   6������o�   ��� 7�����o����� ��Ȁ� �
   |�Ȁ� ���   7�����o�   ����������w���� ��$�   	?�   |�$�   	?���  �������t   ��������������� _@$�   	?�    @$�   	?���   ��������   ��������������@�@$�   	?��    @$�   	?���  ��������   ����ݿ���������@�A@"@   ?�� �@"@   ?��?�  �ݿ������   ��������������_ A@r@ � �> ��@r@ � ���  ��������   ��������ݠ���� @��  � "_�����#�  � "_��    \�����ݠ   ���������|����  ��    $��  ���?�    $���     @������|  ��������������  ��    D�h  ���?�    D�g�     @�������  ?���w����v������ "_��    � R   �����    � M�      w����v��  ?��������n����� _�H    ��W@  ����H    ��J�     �����n�  ?������������� O�$   #��@  ����$   #���     0������`  ?���~����������/�"   '�@@ ����"   '�     ~������@  �������������8'�  G� ��@����  G� @   ������ @8����w����p ������@  ��@�@@����@  ��?      �w����p �  8����9���������� 2�0  c�A  @����0  c�>      �9������  8�������{������ �� �#��  ����2� �#�  @   ����{�   8?����|?�������� ���@�
  ��������@�  p0  �|?���   ����@�������� ��`?�1�y  ������`?�1�x   x�  @����    ��������<����  � ��2������ ��0  ��  ����<�    �����>|������  !����`��������� ��   �>|���    �����~������  ������7�(�� ?���7� ���   @~���    �������<���� � D��  ��I��� ;�  ��@��|   `���<�    ����� �|��� � .O��������� ��������~  0� �|a    ������ > ���� � $&����!  ���� ����� ��~   �� > �    ��������?����@� �~���@ o�@  ��~�� ?���   ���?    �����p��?����A� ��~���� �A  ���~�� ���   p��?    ������������#� o�~�rA  �#� �o�~�q������   ����   `?�����?����0�� �����"  #ȟ� ����������`    `�0   0`?����������0�� W���0  ȟ�  ����/�����`    (��   0�����������hO� �1���`�@�O�  ��������   ��  ?h������������hO� ��p��4 ��O�    p��w��� ��    ��    h�������������'� ����B  � '�  ��O����� �    �0�p   ~������� �������#� ����x�  #� � ����� �      �    ������������������  �� @� � p � ��@�      ��    ������������������ ���� �@� �   � �@�            ����������������x�  a0 @�� ���� � ?���           �xw��������������p�x� ��  ��x ���|  ��w�          �p{�������������.��p@    ��p ����    ��{��           .�;���������������  @ � :  ?��  ?���   ��;��           �=�������������=��� �  �� �� � >  ��=��           =��������������}��	  �� @�� � ���  �  � ��           }������������� ��� 8   �� ���� �� @ � ��       @  �����������������    �@� ���� ��  � ��         ������������������    � � ��� ��   � ��         ��p������������』�    � 0x � ���� ��   x �p         ���?���������������_�    @ @p � _��� ���  p ?�         ?������������������?�  @� > � ?��� ���    �         �������������?����� �  �~ � �����  � ��      �?������������������   � � �� ���   �        ���� ��������������`     >� � �� ���  � �      ���~���������������    �� � �� ���?  �~�       ��I� ��������� ����� |    �� �  |� ����   ���       ��� ?�������� �����<�   ��� �  <   �����   ��       �� �������� ����� x   ���?� �   @ ����  �?���      �I� �������������� � � � �   x ���    ���    ���� � ����� ����������� �  ���� �    �    ���� �� ��?�� ���� p��������(�   p�� ��  (m���   ?�����      } }   ������� ���������p�� �   �  �p    ��� ����� � ������ ������~���� �  ��� �   �7� �   ��rI� � ?������ �����ǀ ��� �  ���  �    � 8    ���� � ?������ ������   ���� �  ����  �   �      ��� �������������7��    �?� �  7�?��    �  m��      �͵� ?�������������G�    ��(�  G���  � (���       ���� ~|���������c����    ���0b ����  � 0��|       >��������������#��     3�� " ���  ��  m��       ������������� ��#��  �� "   ��  ��  ���         ������������� ?�#� � ���"   �� ������       ?��<�������������C�   @��B    ��  ?��=o��         ��8�����������/�pG�p    @ �?�F p  ��  ?����9���         /�px?����������7�p���`    � ?��� �  ��  ����y��         7�pt~����������{�8����    � ����  ��  ����u~          {�8��������������8�    �@�
�  ��  �����           ��8��������������� 8   ��� ��  �_����        @ ���������������|�  �� @����  �   ��� ����           |��������������"�� �  @C�"�  �� ��� C���           ?���?������������$?�@ � :   !�$?߀  ����� !���           �������������� H_�    ��H_��   ����� ����            �������������� HO� ��  	��HO� ��?������          oy���������������  a0 @�x����  �����xox            �^��������������� ���� ��8���   �� �8^�            ����������������B  �� �B���  x � ���     ��     ������� ������B @���x� �B�����  |  ���     �    �{������| ������� �σ��B  ����\O���<  {�   @0| p    �w������|������p� �L��q�4 ��������p   �w�   �|�     p������@|������x �1���`����?����   ?���  @|�   x�������|������8  F?��? ?����?��?   ���   9�|��    8�������|�?����  �?��?�"  ?@��?��?�  @��   g�|�0    ��������<������>@ x��?�A   >?��x��?�>   ��  ��<�   ؀�����<�w������ ������ �� ����   �   �<�v   ������<�{������ �����@ h������?� �   �<�{   ������ �������� $'���!  �������� x    � ���  ������������� .I��������	����@ �   6���a  ����� ����?����� D��  ��� ���  ����    n ����0  ����� ��������� ����`�<� � ?  �`�<���     _ ����  ������|�������� !@���` �  @�����     ��|���   ���������=������ @> ��� �  @> ����    �����=�   �������@7����� �`?�1��  ��   �`?�1�����   ���@6   p����|?���{����� ����
  ��  �������8   �|?���z   @��������{������8 ��! �?�  �0 �! �?@��x�  ����{��    ��������������� 3�F0  cA  x  ��F0  c ����  ��������   ���� w����w�������@  �@�@x  ���@  � ���   w����w��   ���� ���������8'�� D ��x ��� D _��  ������ @ ���� ���������� (�" �$�@@8  ��" �$�?���   �������@   ����������݀���  H~$ �"�@ 8  �~$ �"�?���  7������݀`   ���������n ?���  PH   ���@ 8  
�H   ���?��� /�����n "   �����w����v ?���  "P�   ���  8  ��   ������  /�w����v     ����������� ���@  �	   D��     	   D����  _�������    ����������� _���@  �	    $��    <	    $����  C������� P   ���m�����݃����� @��  "|(�� ??�  "| �   @m�����݃�   �������������� A�@ `>� >�@ `�    ��������  �����z����������A�@ �  �� >�@ �        ���������  ���������������� A 	 � ��� G 	       ��������  ���������ߏ���� _� !  	 v ��� '  	 q�     ������߈   ��� ��������� ��� @ 	/� � �� @ 	/��     ������   ���|7�����`���� ��Ȁ���� � �Ȁ�����    |7�����`   �����` ��`���� ��I������ � �I�������    �������`   �����?���`���� ��I���� � �I�������    �������`   �����  @�`���� ��I���� � �I�������    �������`   �����?���`�������I ����H �I �����    �������`   ��� 6���?��`��������  @ ���~���  � ��P  � 6������`@ ��� 6���_��o���������  )  �
H ��  '� �	�     6������o�   ��� 6���o��o����� ���  I� �
 � ��  W� �	�     6������o�   ��� 6��zw��o����� ���  �� �
 � ��  �� �	�     6������o�   ��� 6�����o����� ��� 	� �
 � �� � �	�     6������o�   ��� 7�����o����� ��Ȁ� �
 � �Ȁ� �	�     7�����o�   ����������w���� ��$�   	?� � �$�   	?��    �������t   ��������������� _@$�   	?� ��@$�   	?��     ��������   ��������������@�@$�   	?�� ?�@$�   	?�  �  ��������   ����ݿ���������@�A@"@   ?��? >@"@   ?�  �  �ݿ������   ��������������_ A@r@ � �>  >@r@ � ���  ��������   ��������ݠ���� @��  � "_��� ?#�  � "_��   \�����ݠ   ���������|����  ��    $��  � ?�    $����   @������|  ��������������  ��    D�h  � ?�    D�`��   @�������  ?���w����v������ "_��    � R   � ���    � @��    w����v��  ?��������n����� _�H    ��W@  � 
��H    ��B?��   �����n�  ?������������� O�$   #��@  � ��$   #��?��   0������`  ?���~����������/�"   '�@@ � ρ"   '��?��   ~������@  �������������8'�  G� ��@���  G� _�  ������ @8����w����p ������@  ��@�@@� ��@  �� ��   �w����p �  8����9���������� 2�0  c�A  @� ��0  c� ���   �9������  8�������{������ �� �#��  �� � �#�@��@   ����{�   8?����|?�������� ���@�
  ��  ���@����p0  �|?���   ����@�������� ��`?�1�y  �    ��`?�1�x���x�  @����    ��������<����  � ��2��   � ��1����  ����<�    �����>|������  !����`�   ��������   �>|���    �����~������  ������7�(�  ? ?���7�'����   @~���    �������<���� � D��  ��I�� ���  ��F���|   `���<�    ����� �|��� � .O���������������@ ��~  0� �|a    ������ > ���� � $&����!  ���������� {�~   �� > �    ��������?����@� �~���@ o�@���~��?� �   ���?    �����p��?����A� ��~���� �A�� ��~��  �   p��?    ������������#� o�~�rA  �#���o�~�p>  ��   ����   `?�����?����0�� �����"  #ȟ�������  �`    `�0   0`?����������0�� W���0  ȟ�������    �`    (��   0�����������hO� �1���`�@�O���?����    ��   ��  ?h������������hO� ��p��4 ��O���pp��    ��    ��    h�������������'� ����B  � '����O��<   �    �0�p   ~������� �������#� ����x�  #�����  |   �      �    ������������������  �� @����  x �  @�      ��    ������������������ ���� �@���   ��  @�            ����������������x�  a0 @����  ������           �xw��������������p�x� ��  ��x� ��?���w�          �p{�������������.��p@    ��p?�   ������{��           .�;���������������  @ � :  ?�� �  ������;��           �=�������������=��� �  ��  �� ���?�=��           =��������������}��	  �� @�� �  �   ���� ��           }������������� ��� 8   �� �  ��  �_�� ��       @  �����������������    �@� �  ��  ��� ��         ������������������    � � �  ��  ��� ��         ��p������������』�    � 0x � �� ��  ��x �p         ���?���������������_�    @ @p � _� ��  ?��p ?�         ?������������������?�  @� > � ?� ��  ?�   �         �������������?����� �  �~ � � �� � � ��      �?������������������   � � � ��  �  �        ���� ��������������`     >� � � ��  �  � �      ���~���������������    �� � � ��  ?  �~�       ��I� ��������� ����� |    �� �  | ��  �   ���       ��� ?�������� �����<�   ��� �  < ?��  ��   ��       �� �������� ����� x   ���?� �   G��  ��  �?���      �I� �������������� � � � �   x�  �    ���    ���� � ����� ����������� �  ����  �    �    ���� �� ��?�� ���� p��������(�   p�� ��  (m���   ?�����                                                                                                                                          