��j  �V�                                x                                                                       x                                                                       x                                                                       x                                                                      � � 0                                                                 � � 0                                                                � � 0                                                                  � � 0                                                                 � � 0                                                                � � 0                                                                � � 0                                                                 � � 0                                    0                        /    ��<y��;�Ǚ�                              /                            ��<y��;�Ǚ�                              8                        '    ��<y��;�Ǚ�                                                           ��<y��;�Ǚ�                                                      o�   y�f̀3m�l�6      /                        o�                           y�f̀3m�l�6      .                        0�                       O    y�f̀3m�l�6      �                       _                             y�f̀3m�l�6                               @                       _�   �~���3m��6      �                       _�                            �~���3m��6      X�                       a�                       @   �~���3m��6      ?                        >                             �~���3m��6                              ��                       ��                       \                        ��                       @                        ^                        �                       ��   �`���33m��6      9�                       \                                                                         @                       ��                       ��                      ��                       @                        ��                       �`                      <�   ͛f́�33m�l�6      v`                      |�                                                0                        ��                      x                       k�                      x                       ��                      c�                      ��                       y`   x�<x��3m�Ǚ�m�    ��                       ��                                                a�                      �                      ��                      q�                      ��                       `                      {�                      ��                      s�                       �f                      p`                                                ``                      �                      ��                     �~                      ��                                            ��                      ��                     ��                      ��                     �                                                �                      �                     ���                     ���                     ���                                            ��                     �                     ���                     �`                     �                                               �                      ��                     ��x                     ���                     ��x                      �                     ��                     ?��                     	��`                     ��                     �a�                                              ��                     ��                     ���                     ���                     ��                       `                     �g�                     7��                     ���                     a�f                     �`                                                `                     ��                     ���                    ��~                     ���                                           ?��                     ���                    ���                     �`�                    �                                                                     0?��                    /����                    ?���                    /����                                           ���                    8���                    '?���                    @`                     �                                                                     ��                    o���x                    /_���                    o���x                      �                    ._���                    0���                    O?��`                    � �                    _ a�                                               �                     g�g�                    _���                    �y�                    _���                        `                    X�g�                    a��g�                    g��                    ?  f                    >  `                                                `                    @� �                    ?� �                   \W ~                    ?� �                   @@                      ^_ �                    c� ��                   � �                    9�  �                   \D                                              @                       { �                   � ��                   7 ��                   � ��                                           9; �                   { �                   � ��                   �  `                   � �                                                                    = ��                   � �x                   � ��                   � �x                      �                   
= ��                   } ��                   	� �`                   P  �                   �  a�                                               �                   �  g�                   �  �                   �  y�                   �  �                       `                   �  g�                   �  g�                   �  �                    P   f                      `                                                `                    ^� �                    w� �                   ]� ~                    w� �                                          ^� �                    ~� ��                   W� �                    (   �                   	                                                                      � �                   7� ��                   � ��                   7� ��                                          � �                   >� �                   � ��                   (   `                   	  �                                                                    @ ��                   � �x                   � ��                   � �x                      �                   @ ��                   @ ��                   � �`                      �                   �  a�                                               �                   @  g�                   �  �                   �  y�                   �  �                       `                   @  g�                   @  g�                   �  �                       f                   �  `                                                `                   �  �                   �  �                  `  ~                   �  �                                         �  �                   �  ��                  �  �                   
    �                  @                                                                     �  �                  �  ��                  `  ��                  �  ��                                         �  �                  �  �                  �  ��                  
    `                  @  �                                                                   �  ��                  �  �x                  �  ��                  �  �x                      �                  �  ��                  �  ��                  �  �`                      �                      a�                                               �                  �   g�                  �   �                  �   y�                  �   �                       `                  �   g�                  �   g�                  �   �                       f                      `                                                `                  �  ��                  �����                 �   ~                  �����                  �                      �  ��                  �������                 x  ��                  ���� �                  �                                               �                      �����                 ������                 �������                 ������                  �                      �����                 �����                 ������                 �    `                  �  ��                                            �                       ���� ��                 �  ��x                  �������                 �  ��x                  _��� �                  ���� ��                 ���� ��                  �  ��`                 _��� �                  _����a�                                           _��� �                  ���� '�                 �������                  �������                 �������                  @     `                  ���� '�                 ���� '�                  �������                 @     f                  @  ��`                                           @     `                  ��� 	�                  �������                 `  ��~                  �������                                         ��� 	�                  ���� 	��                 _������                  �     �                    ��                                                                   p                      ��������                 �������                 ��������                                         p    �                 �    �                 _������                  �     `                 /������                                                                   ?�������                 o������x                 ?��� ��                 o������x                      �                 ?�������                 �������                 /������@                 P     �                      a�                                               �                 =     g�                 o     �                 ;     y�                 o     �                       `                 =     g�                 }     g�                 /     �                 P      f                      `                                                `                 �    �                 7�    �                �    ~                 7�    �                                       �    �                 >�    ��                �    �                 (      �                	                                                                      �                     7�    ��                �    ��                7�    ��                                       �    �                >�    �                �    �                 (      `                	     �                                                                 @    ��                �    �x                �     ��                �    �x                      �                @    ��                @    ��                �    �@                      �                �     a�                                               �                @     ��                �    ��                �    y�                �    ��                      @`                @    ��                @     ��                �    ��                       f                �    X`                                                `                �     ��                �     ��               `     �~                �     ��                     @                �    Y�                �     ���               �     ��                
      ��               @     F                                               @                �     .�               �     ���               `     ǟ�               �     ���                                      �     N�               �     ~�               �     ���               
      �`               @     ��                                               @                �     )��               �     ]�x               �     a��               �     ]�x                      �               �     ���               �     y��               �     �`                     p�                     $a�                                               �               �     Pg�               �     l�               �     `y�               �     l�                      `               �     ���               �     xg�               �     D�                     x f                     `                                                `               �     �               x     l?�              �     0~               x     l?�               �                     �     T�               �     <��              x     @7�               �     8 �               �     P&                                         �                     �     (
�              x     67��              �     0��              x     67��               �                    �     P�              �     <�              x     "#��              �     <`               �     
)�                                         �                     �     	��              �     67�x               �     ��              �     67�x               @     �               �     *+��              �     ��               �     "#�`              @     �               H     **a�                                        @     �               �     g�              �     l�               �     y�              �     l�               @      `               �     (
g�              �     8g�               �     D�              @     < f               H     T`                                        @      `               z     �               �     l�              v     ~               �     l�                                    z     T�               �     8��              ^     D�               �     8 �              $     T                                                              z      �              �     ���              v     ��              �     ���                                     z     �              �     p�              ^      ���              �     x `              $     ��                                                              =     
 ��              o     ��x              ;     0��              o     ��x                     �              =     
���              }     ���              /     �`              P     p �                   ( a�                                              �              =     @ g�              o     � �              ;     0 y�              o     � �                   @  `              =     
( g�              }     � g�              /      �              P     �  f                   P `                                               `              �    @ �              7�    � �             �    ` ~              7�    � �                  @                �    P �              >�    � ��             �     �              (     �  �             	     P                                             @                �    � �             7�    ` ��             �    ` ��             7�    ` ��                   �                �    P �             >�    � �             �      ��             (     �  `             	      � �                                            @                @       ��             �    � �x             �    � ��             �    � �x                      �             @    � ��             @    � ��             �      �`                  �  �             �       a�                                            �  �             @        g�             �        �             �     �  y�             �        �                       `             @    `  g�             @        g�             �        �                   �   f             �        `                                                `             �        �             �        �            `        ~             �        �                                   �    �  �             �        ��            �        �             
          �            @                                                                     �        �            �        ��            `        ��            �        ��                                   �        �            �        �            �        ��            
          `            @        �                                                             �        ��            �        �x            �        ��            �        �x                      �            �        ��            �        ��            �        �`                      �                      a�                                               �            �         g�            �         �            �         y�            �         �                       `            �         g�            �         g�            �         �                       f                      `                                                `            �         �            x         �           �         ~            x         �            �                      �         �            �         ��           x         �            �          �            �                                               �                      �         �           x         ��           �         ��           x         ��            �                      �         �           �         �           x         ��           �          `            �         �                                      �                       �         ��           �         �x            �         ��           �         �x            @          �            �         ��           �         ��            �         �`           @          �            H          a�                                     @          �            �          g�           �          �            �          y�           �          �            @           `            �          g�           �          g�            �          �           @           f            H          `                                     @           `            z          �            �          �           v          ~            �          �                                   z          �            �          ��           ^          �            �           �           $                                                                       z          �           �          ��           v          ��           �          ��                                   z          �           �          �           ^          ��           �           `           $          �                                                             =          ��           o          �x           ;          ��           o          �x                      �           =          ��           }          ��           /          �`           P           �                      a�                                               �           =           g�           o           �           ;           y�           o           �                       `           =           g�           }           g�           /           �           P            f                      `                                                `           �          �           7�          �          �          |           7�          �                                 �          �           >�          ��          �          �           (            �          	                                                                      �          |           7�          ��          �          �           7�          ��                                 �          �          >�          �          �          �           (                       	           �                                                           @          ��          �          ��          �          ��          �          ��                                  @          �          @          ��          �          ��                      �          �           `                                                            @           g�          �           �          �           w�          �           �                                  @           h          @           o�          �           w�                      �          �                                                                       �           �          �           ��         `           �          �           ��                                 �                     �           ��         �           �          
            ��         @                                                                        �           ��         �           ��         `           ��         �           ��                                �           �         �           ��         �           ��         
            �`         @                                                                      �           ��         �           �x         �           ��         �           �x                      �         �           �         �           ��         �           �`                     ��                      �                                               �         �           ��         �           ��         �           ��         �           ��                       `         �           �         �           ��         �           ��                     �f                       `                                                `         �           ��         x           ?��        �           �~         x           ?��         �                      �           0�         �           ?���        x           ��         �           ��         �                                               �                      �           ��        x           ?���        �           ���        x           ?���         �                      �           (�        �           ?��        x           ���        �           �`         �            �                                   �                       �           ��        �           ?��x         �           ���        �           ?��x         @             �         �           $��        �           ?��         �           ��`        @           ��         H             a�                                  @             �         �           < g�        �           ��         �           < y�        �           ��         @              `         �           C�g�        �           �g�         �           < �        @           <  f         H             `                                  @              `         z           < �         �           ~ �        v           < ~         �           ~ �                                z           B �         �           ~ ��        ^           < �         �           <  �        $                                                                       z           < �        �           ~ ��        v           < ��        �           ~ ��                                z           B �        �           ~ �        ^           < ��        �           <  `        $             �                                                          =           x ��        o           � �x        ;           x ��        o           � �x                      �        =           � ��        }           � ��        /           x �`        P           x  �                      a�                                               �        =           x  g�        o           �  �        ;           x  y�        o           �  �                       `        =           �  g�        }           �  g�        /           x  �        P           x   f                      `                                                `        �          x  �        7�          �  �       �          x  ~        7�          �  �                              �          �  �        >�          �  ��       �          x  �        (           x   �       	                                                                      �          �  �       7�         �  ��       �          �  ��       7�         �  ��                              �           �       >�         �  �       �          �  ��       (           �   `       	              �                                                        @          �  ��       �         �  �x       �          �  ��       �         �  �x                      �       @           ��       @         �  ��       �          �  �`                  �   �       �              a�                                               �       @          �   g�       �         �   �       �          �   y�       �         �   �                       `       @            g�       @         �   g�       �          �   �                  �    f       �              `                                                `       �          �   �       �         �   �      `          �   ~       �         �   �                             �            �       �         �   ��      �          �   �       
           �    �      @                                                                     �              �      �         �   ��      `              ��      �         �   ��                             �         �   �      �         �   �      �              ��      
                `      @              �                                                       �             ��      �            �x      �             ��      �         �   �x                 �    �      �         �   ��      �            ��      �             �`                     �                      a�                                               �      �               g�      �             �      �               y�      �         �    �                �     `      �         �    g�      �             g�      �               �                       f                      `                                                `      �               �      x             �     �               ~      x             �      �                    �             �      �         �    ��     x          �    �      �          �     �      �                                               �                      �          �    �     x         �    ��     �          �    ��     x         �    ��      �         �           �         �    �     �         	    �     x             ��     �              `      �               �                                �                       �          �    ��     �         �    �       �          �    ��     �         �    �       @         �     �      �         �    ��     �         	    ��      �             �      @              �      H                �                               @                �      �          �     A�     �         �     �      �          �     A�     �         �     ~<      @         �             �         �     @      �         	     �      �              A�     @              ?�      H                                                 @                        z                �      �              ?�      v                �      �              =�                     �      z              �      �         �     ?�      ^          �     �      �          �     ?�      $                �                       �                       �      z                0      �              ><      v                0      �         �     :,                �            z         �            �              ?�      ^                �      �                ?�      $                                                                       =               �      o              >�      ;               �      o         �     :,                �            =         �            }              ?�      /               �      P               ?�                                                                            =                0      o         �    �<                      0      o         �    �,                             ?         �            }         �    ��      /                �      P               ��                                                                            �        �    ��      ?�        �    ��               �    ��      ?�        �    ��                       �      �            ��      >�        �    ��      �        �    ��      .         �    ?�                      �                       �                       �       �        �    ��      ?�        �    ~?�                �    ��      ?�        �    ~><                      �        �            �       ?�        �    ��       �        �    �      ?         �    q��                      �                                                �       @        �    �       �        �   ���      �        �    �       �        �   ���                              �            �       @        �   ���      �        �    q�                �   ��      �                                                                                 �   ��       �        �   ��       @        �   �?       �        �   ��                       p        @           ��       �        �   ��       @        �   ��       �        �   p        @              p8                                                p                  �   �8       �        �   ��                 �   ��       �        �   ��                      �                     �8       �        �   ��8                 �   �       �        �   �                       ��                                               �                  �   ���       �        �  ���                �   ���       �        �  ���                                0           ���       �        �  ���        0        �   ���       �        �                                                                                            �  ��        �        �  ?�        �         �  �~        �        �  ?�                       �         �          ��        p        �  ?��        �         �  �        `         �  8�         �             �p                                                �                   �  ?�p        �        � ���        @         �  ?��        �        � ���                                H          ?�p        �        � ��p        H         �  8��        �         � �          @            �                                                                  � ��        �        � ���        �         � ��        �        � ���                      8          
�         ��        \        � ��        �         � ���        X         � 8          
�            8                                                8          �         � �         �        � ~?�         �         � ��         ~        � ~?�                      �          &         �         �        � �         �         � ?�         �         � q�          $           ��                                               �                   � ��         �        ����         �         � ��         �        ����                                 
�         ��         Y        ����         �         � q��         X         ��           
�                                                                       @      `���          ��   ��!����          D�      @��?          ��   ��!����                   @  p           G�      a ���          �@   ��a����          G�       ���          �    ��@�p           D�      @  p8                                            @  p            �    �� ?��8          ��   �������          �`        ?���          ��   �������                     �           ��    �� �_�8          �   �������8          ��    �� ?��          ~    � �?��           �@         ��                                              �            �   � ����          ��   � �����          8        ߏ�          ��   � �����                                 �   � ��?��          ��   � �����          �   � ����          �         �            "                                                                    ��      ߎ           �?�����������           �      �~           �?�����������             �                    ��      �?�           �������������           �>        ��            	����������            �          p                                      �                       ����������p            ������������            
y����������            ������������             <                       ����������<p            �����������p            �����������             <      �             
=         �                                      8                       {��������À            �      ���            ���������߀            �      ���             ��������               ����������#�            ����������            �      ߀             ���������             ���������                                      ��������               ����������             �����������              q���������             �����������                                      ����������<             �����������             ����������                     �              p                                                                          1����������              ����������              ~        ?�              ����������                                       q���������`              1����������              ����������                     ?�              N                                                                                                 ����������              ���������               ����������                                            �                      ?�              ���������                                       ���������                                                                 ���������               ���������               ���������               ���������                                      ���������               ���������               ���������                                                                                                                  ?�    `                  ?�    `                  ?�    `                  �����                  �����                  �����                  ;�                       ;�                       ;�                                                                                                  ?������                  ?������                  ?������                                                                                             ?������                  ?������                  ?������                                                                                             �    x                  �    x                  �    x                                                                                          �    h                  �    h                  �    h                                                                                                   <                        <                        <                                                                                                4                        4                        4                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �0�߀                     ���                   �o��7�                                                                                                                                                                                                                                                 �0��                      ��                    llll6                                                                                                                                                                                                                                                  �x��                      �                    llnv                                                                                                                                                                                                                                                  �x��                      �                    llnv                                                                                                                                                                                                                                                  ����                      ��                    ��o��                                                                                                                                                                                                                                                 ����                      ��                    llo�                                                                                                                                                                                                                                                  ����                      ��                    llm�                                                                                                                                                                                                                                                  ����                      �0�ـ                   lllm�                                                                                                                                                                                                                                                  ����                      ��Ϙ�                   �lg�7�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        
 �       �              T                   T            
                                                                                                                                                                                                                                         �       �              $                   $            
                                                                                                                                                                                                                                        
       �              ""                   ""            
                                                                                                                                                                                                                                        *,rǜ���q�          ""T��+��$�y���       ""T��+�3�� �<�zq�                                                                                                                                                                                                                                      *�(����R�           ""T) ��((�"�)�       ""T) ��,�RQ �D��R                                                                                                                                                                                                                                      �*"z(�"����           !TT�'��)�0>���       !TT�'���R_ �D��                                                                                                                                                                                                                                      �*"�(�"��D�           !TT	(��*(( �)       !TT	(���RP �E���                                                                                                                                                                                                                                      D*��(����R�            �T)(��*(�"�)�        �T)(��(�RQ �E��R                                                                                                                                                                                                                                      D*"z'�����q�           �T�'����"Ay���        �T�'��ȣ�N �<�zq�                                                                                                                                                                                                                                            �                             �                        @                                                                                                                                                                                                                                                                               �                        x                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             @                     @                                                                                                                                                                                                                                                        �                    @                     @                                                                                                                                                                                                                                                        �                    @                     @                                                                                                                                                                                                                                                �㓘�v8�               �99��X�c�              �99��X�c�                                                                                                                                                                                                                                             ATP%QID�               (EEQe�H              (EEQe�H                                                                                                                                                                                                                                             ATP_I|�               (EEE���              (EEE���                                                                                                                                                                                                                                             ATP	PI@�               (EE �E�              (EE �E�                                                                                                                                                                                                                                             ATP%QID�               (EEQE�H              (EEQE�H                                                                                                                                                                                                                                              �@㓐�NI8�               �99�D䓈              �99�D䓈                                                                                                                                                                                                                                                        �                                                                                                                                                                                                                                                                                                                                                                                                                                           