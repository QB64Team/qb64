��]  ԶT�                            �    �   0   0 �                                                       �    �   0   0 �                                                       �    �   0   0 �                                                       �    �   0   0 �                                                       `  � �0   0 �                                                       `  � �0   0 �                                                       `  � �0   0 �                                                       `  � �0   0 �                                                          � �0   0 �                                                          � �0   0 �                                                          � �0   0 �                                                          � �0   0 �                                                       �����;`9ͳ�y��<y�p                                                      �����;`9ͳ�y��<y�p                                                      �����;`9ͳ�y��<y�p                                                      �����;`9ͳ�y��<y�p                                                      ��6l ����m��`�0fͳ`                                                      ��6l ����m��`�0fͳ`                                                      ��6l ����m��`�0fͳ`                                                      ��6l ����m��`�0fͳ`                                                                                                                                                                                                             o������1���}�0`ͳ`                                                                                                                                                                                                                                                                                        l������ ͛0`ͳ`                                                                                                                                                                                                                                                                                       l�6l���`m�6`͛0fͳ`                                                                                                                                                                                                                                                                                       Ǚ����308�3�}��<y�f�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     �                                                                         �                                                                         �                                                                         �                                                                        �                                                                        �                                                                        �                                                                        �                                                                        �                                                                        �                                                                        �                                                                        �                                                                                                                    @                                                                     @                          �           ?                               @                                                                      @                          2�         >(                   
            �           
               5�         >(                   
            �           
               7�         n8                               �                          2�         .(                   
            �           
               =@         �D                                                        {@         �D                                                        �         �|                              �                          @         �D                                                       >
�         �                  *          �          *              �
�         Ш                  *          �          *              �         ��                  6          `          6              
�         ��                  *          �          *               �          �                  (D          �@          (D              ~          �                  8D          �@          8D                          ��                  (|          ��          (|                          �                  (D          �@          (D              2          G�                   d�          L�          d�              �2          K�                   |�          ̀          |�              .          @��                  D�          K�          D�              "          @�                   D�          H�          D�              �          '�@                  cP          5           cP              ��          e�@                  ?P          �           ?P               ��          ��                  C�          ;           C�               O�          �@                             1                         ��         ��                  ��          
           ��              o�         ,��                  ��          	�           ��              ��         ��                  �          :           c�              ��         ��                  �                      �              	Op          ��                  p�                    p�              ��         �                  ��          �          l�              �p          4w                  ��          <           ��              p          w                   `�                     `�              B�0         <s                  �@          /�          �@              M��         �?                  4@          -D          �@              G�0         h�                  ��          �          ��              B0          3                   �@                     �@              %+8         z�                 �           ^B          �               kq�         n߀                 x           Z          �                         �р                 ��          =�          ��              	          @р                 �                     �              8         ��                 B@          �$          �@             7,�         �߀                 �@          �          @@             <         ���                 s�          {<          ��                      ���                 �@          0           @              ��0         	��                  ��         x          ��             ��p         ��                  ��         h          ��              <~          G@                  �          �          a�                                             �          `           �             ,T          CǢ                  -           �           /               ܼ          KGb                  3�          �           -               x�          F��                  =�          �           �               @          B                               �                          R�          '�@                  Z           �           ^               �x          f��                  g�          �           Z                ��                             {�          �           =�               @�                                        �                          �P         �                  �           �           �               r�         -�                  �           @           �               ��         :                   �           �           {               �                             8                       0               	J�          ��                  h           �          x               ��         ��                  �           �          h               ��          4t                  �           `           �                          0                   p                       `               B�@         <z                  �           /           �               M��         �v                  <           -           �               G��         h�                  �           �          �               B           `                   �                       �               %*�         z�                  �           ^           �               kw�         n�                  x           Z           �               �          ��                  �           =�          �                          @�                  �                      �                        ��                  @           �           �              7/          ��                  �           �           @              ?          ��                  p           {           �                        ��                  �           0                          ��          ��                  �          x           �              ��          ��                  �          h           �              �~          G@                  �           �           `              �                                          `                           �T          Ǡ                  m           �           o                ܼ          G`                  s�          �           m               ��          >��                  }�          �           ^�               �@                             N           �           L                r�          �@                  �           �           �                wx          ��                  �          �           �               ��                             ��          �           ��               `�                             �           �           �               1P          C�                 �           �          �                2�          �                 �           @          �               ��          ?:                  �           �          �                1                             �                      �               :�          #�                  �           �          �                =�          �                   �           �           �               ��          �                   �           �           �                :           �                   �           �           �               =@          3�                  �           (�          �               ?�          #�                  |           '�          |               ��          o�                             @                         <           #�                               @                          ��          {�                  �           \�          �               ?�          c�                  >           [�          �               w�          �p                  �           8           �               6           C`                  �                      �               
           ��                  o           ��          �               ?           ��                  �           ��          _               3          �0                  A           x          �               3           �0                  �           0                         ?�         ��                  ��         y�          ��              ,_�         ��                  �         h�          ��              <Q�         E                  �          �          a�              �                            �          `           �              (_�         ��                  -          ��          /               X��         F�                  3�          �p          -               x��         �                  =�          �          �                @�                                      �                         P�@         �t                  Z          �`          ^               ��         ��                  g�          �           Z               ��@                           {�          �           =�               @�@                                     �                          �S          �                  �           �           �               b�         �                  �           @           �               ��          :                   �           �           {                �                              8                       0               B�          =                 h           �          x               ��          ;                 �           �          h               ��          4t                  �           `           �                          0                   p                       `               �@          <z                  �           /           �               ��          4v                  <           -           �               ��          h�                  �           �          �                           `                   �                       �               
�          x�                  �           ^           �               �          h�                  x           Z           �               �          ��                  �           =�          �                          @�                  �                      �               
           ��                  @           �           �               /           ��                  �           �           @               ?          ��                  p           {           �                          ��                  �           0                           *          ��                  �          x           �               ,^          ��                  �          h           �               <~          G@                  �           �           `                                                         `                           (T          Ǡ                  -           �           /                X�          G`                  3�          �           -                x�          ��                  =�          �           �                @                                         �                           P�          �@                  Z           �           ^                �x          ��                  g�          �           Z                ��                             {�          �           =�               @�                                        �                           �P          �                  �           �           �               b�          �                  �           @           �               ��          :                   �           �           {                �                              8                       0               B�          =                  h           �          x               ��          ;                  �           �          h               ��          4t                  �           `           �                          0                   p                       `               �@          <z                  �           /           �               ��          4v                  <           -           �               ��          h�                  �           �          �                           `                   �                       �               
�          x�                  �           ^           �               �          h�                  x           Z           �               �          ��                  �           =�          �                          @�                  �                      �               
           ��                  @           �           �               /           ��                  �           �           @               ?          ��                  p           {           �                          ��                  �           0                           *          ��                  �          x           �               ,^          ��                  �          h           �               <~          G@                  �           �           `                                                         `                           (T          Ǡ                  -           �           /                X�          G`                  3�          �           -                x�          ��                  =�          �           �                @                                         �                           P�          �@                  Z           �           ^                �x          ��                  g�          �           Z                ��                             {�          �           =�               @�                                        �                           �P          �                  �           �           �               b�          �                  �           @           �               ��          :                   �           �           {                �                              8                       0               B�          =                  h           �          x               ��          ;                  �           �          h               ��          4t                  �           `           �                          0                   p                       `               �@          <z                  �           /           �               ��          4v                  <           -           �               ��          h�                  �           �          �                           `                   �                       �               
�          x�                  �           ^           �               �          h�                  x           Z           �               �          ��                  �           =�          �                          @�                  �                      �               
           ��                  @           �           �               /           ��                  �           �           @               ?          ��                  p           {           �                          ��                  �           0                           *          ��                  �          x           �               ,^          ��                  �          h           �               <~          G@                  �           �           `                                                         `                           (T          Ǡ                  -           �           /                X�          G`                  3�          �           -                x�          ��                  =�          �           �                @                                         �                           P�          �@                  Z           �           ^                �x          ��                  g�          �           Z                ��                             {�          �           =�               @�                                        �                           �P          �                  �           �           �               b�          �                  �           @           �               ��          :                   �           �           {                �                              8                       0               B�          =                  h           �          x               ��          ;                  �           �          h               ��          4t                  �           `           �                          0                   p                       `               �@          <z                  �           /           �               ��          4v                  <           -           �               ��          h�                  �           �          �                           `                   �                       �               
�          x�                  �          ^           �               �          h�                  x          Z           �               �          ��                  �          =�          �                          @�                  �                     �               
           ��                  +@          �           +�               /           ��                  ,�          �           +@               ?          ��                  ?p          �           ?�                          ��                  +�          �           +                *          ��                  ^�          �           _�               ,^          ��                  ]�          �           ^�               <~          G@                  ~�          �           `                                             _           �           ^                (T          Ǡ                  �           �           �                X�          G`                  ��          �           �                x�          ��                  ��          �           ��                @                             �           �           �                P�          �@                            �                          �x          ��                 �          �                          ��                            ��          �          ��               @�                                       �                          �P          �                  ��          �           ��              b�          �                  ��          �           ��              ��          :                  ��          �          ��               �                              ��          �           ��              B�          =                  ��          �          ��              ��          ;                   ��          �           ��              ��          4t                  ��          �          ��                         0                   ��          �           ��              �@          <z                  ��          +          ��              ��          4v                  7�          3x          7�              ��          h�                  ��          ?�          ��                          `                   1�                     1�              
�          x�                  �           ^0          �               �          h�                             `�          �               �          ��                  �           }0          �                          @�                  �           0          �               
           ��                  �           �`          �               /           ��                  ^           ��          �               ?          ��                  �           �`          �                          ��                  �           8`          �               *          ��                  T          u@          t               ,^          ��                  �          ��          L               <~          G@                  �          �@          �                                             $           r@                         (T          Ǡ                  .�          �           .�               X�          G`                  1�                     .�               x�          ��                  ?�          �           `                @                             @           �                           P�          �@                  ]           �           ]�               �x          ��                  c�          <           ]                ��                             @          �           >�               @�                             �          �                           �P          �                  �           �           �               b�          �                  ǀ          x           �               ��          :                   ��          �           }�               �                              9           �           8               B�          =                  t           @          v               ��          ;                  �           �          t               ��          4t                  �           �           �                          0                   r                       p               �@          <z                  �           .�          �               ��          4v                             1�          �               ��          h�                  �           ?�          �                           `                   �           @           �               
�          x�                  �           ]           �               �          h�                  <           c�          �               �          ��                  �           @          �                          @�                  �           �          �               
           ��                  �           �           �               /           ��                  x           ǀ          �               ?          ��                  �           ��          �                          ��                  �           9           �               *          ��                  @          t           `               ,^          ��                  �          �           @               <~          G@                  �          �           �                                                         r                           (T          Ǡ                  .�          �           .�               X�          G`                  1�                     .�               x�          ��                  ?�          �           `                @                             @           �                           P�          �@                  ]           �           ]�               �x          ��                  c�          <           ]                ��                             @          �           >�               @�                             �          �                           �P          �                  �           �           �               b�          �                  ǀ          x           �               ��          :                   ��          �           }�               �                              9           �           8               B�          =                  t           @          v               ��          ;                  �           �          t               ��          4t                  �           �           �                          0                   r                       p               �@          <z                  �           .�          �               ��          4v                             1�          �               ��          h�                  �           ?�          �                           `                   �           @           �               
�          x�                  �           ]           �               �          h�                  <           c�          �               �          ��                  �           @          �                          @�                  �           �          �               
           ��                  �           �           �               /           ��                  x           ǀ          �               ?          ��                  �           ��          �                          ��                  �           9           �               *          ��                  @          t           `               ,^          ��                  �          �           @               <~          G@                  �          �           �                                                         r                           (T          Ǡ                  .�          �           .�               X�          G`                  1�                     .�               x�          ��                  ?�          �           `                @                             @           �                           P�          �@                  ]           �           ]�               �x          ��                  c�          <           ]                ��                             @          �           >�               @�                             �          �                           �P          �                  �           �           �               b�          �                  ǀ          x           �               ��          :                   ��          �           }�               �                              9           �           8               B�          =                  t           @          v               ��          ;                  �           �          t               ��          4t                  �           �           �                          0                   r                       p               �@          <z                  �           .�          �               ��          4v                             1�          �               ��          h�                  �           ?�          �                           `                   �           @           �               
�          x�                  �           ]           �               �          h�                  <           c�          �               �          ��                  �           @          �                          @�                  �           �          �               
           ��                  �           �           �               /           ��                  x           ǀ          �               ?          ��                  �           ��          �                          ��                  �           9           �               *          ��                  @          t           `               ,^          ��                  �          �           @               <~          G@                  �          �           �                                                         r                           (T          Ǡ                  .�          �           .�               X�          G`                  1�                     .�               x�          ��                  ?�          �           `                @                             @           �                           P�          �@                  ]           �           ]�               �x          ��                  c�          <           ]                ��                             @          �           >�               @�                             �          �                          �P          �                  �           �           �               b�          }�                  ǀ          x           �                ��          
:                   ��          �           }�               �                              9           �           8                          �=                  t           @          v               ��          �;                  �           �          t                G�          t                  �           �           �                            0                   r                       p               �@         �z                  �           .�          �               ��         �v                             1�          �               �          p�                  �           ?�          �                          p`                   �           @           �              ��         q��                  �           }           �              ��         w��                  <           s�          �               �          pP                   �           @           �                           p@                   �           �           �              ��          ��h                  �           �           �              ��          ���                  �           ��          �                           p                   h           v�          X                           p                              q                          O�         t��                  �          �           �              ��         ���                  �          �           �               8          p�                  �           �           �               8          p�                  �           �           �              G�         t{�                  ?�          �           ?�              ��         ���                  :�          �           :�               8          p�                  /�          �           �               8          p�                  
�           �           
�              @�         t�                  _�          �           _�              ��         ���                  }�          �           ]�               8          p�                  o�          �           /�               8          p�                  �          �           �              �D          �@                  ?�          �           ?�              ��          ���                  O�          �           ?�                                                w           p           w                                                 7           p           7                8          p�                  7           p           7               �          w��                              �           7                                                 8           �           8                                                 0                       0                                                             �                                                                       �                                                                       �                                                                        @                                                                                                                                                    �                                                                                                                                                 �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ��  �         �        �0   � �   �    ` �  �`     �                                                                                                                                                                                                                                      `    �  �   �    6         0      `    �          `      �                                                                                                                                                                                                                                           �  �                 0      `    �      �    `                                                                                                                                                                                                                                            ��>y���|�   >v����y�x    3�<��>g��   ���Ǐ>o����  g�<y�||9���                                                                                                                                                                                                                                  �ٻf́�v�   3f�6lͶ�    �m�fͻf�۶   �m�lٳnك��  3l�f͛v��6�0                                                                                                                                                                                                                                   lٳf����f�   �f͛�lͶ�    ��0fͳf�6   �����lك��  ?o�`͛f��6��                                                                                                                                                                                                                                   lٳf����f�   �f͛lͶ�    60fͳf�6   ����lكm�  0l`͛f��6�                                                                                                                                                                                                                                   lٳf́��f�   �f͛66lͶ�    �m�fͳf�6   �m�lٳlكm�  3l�f͛f�ٳ6�0                                                                                                                                                                                                                                  ϙ�>y���f`   >f����ly�x    3�<��>�3   ���Ǐ>lσ�  g�<y�f|�����                                                                                                                                                                                                                                               0                   �             0 �         �                                                                                                                                                                                                                                            |          0 �                 � |            0           � �                                                                                 