�h  ��Q Q  g�����0   �    �                         �������   @ ?�                        ����d   ��� �      ?�                 n��?���    ?� D    ��                �������   c���                      ���  <���  H����	     `                 _�t  /�`  �t  0�  �   �             ���   ���  @�  �       0 @            ��   >1��  g   ��    ��    �            �\@  <��  �@  = P   #�  ��              ���  �� ��  �   G  ��            /�a  ?� q    �  ���            [��   @q�� $�   `��    ?�              ��  A ���(	�  A��
 @  ~ 0      @     ��   � w��@"  � p   �  �      �     o� �  ;� �& �  8� 8  �  L       �    _�    7� �lD   6� 8 �             ��@    �� XD    @ 8 �             ��H   ��@�H   �  @0 �             ~     ?��0�   @  �p �  �            @  `&  ���`� p7  �  �p �  �          � ��  �*  ��� �:�    p s�   �           ��  ��  ��� ��� `  p p   �     p   @ ��     ���� ���  �  p p   `           �       ���� �   �  p      `            � H �L�  W� L 泀  X  0 ��  0     �@�   � D���~ _� D�3���X  8 ��  0     ���   � � ���k� F�����l  8  a�       @�  �  ��� P+� ��� X,  >� ���    � � @ � #� � /� #���� ,  ����   � �  � ����  � ���   ������   �� �   �  ��� �, �!�  �=���      |   � ?�~`@�, ?� �y��  ��?�?    >  >   � >�>��, ? ~�0  ��ߟ �    <     � z@�/  Z�\ z�b��[   �^�_ �    x     � ��� 
�\ ��P�    z�� �     �    �  ��  �\      �����         �  ��� �\  X     ����� �          �  s�  �^  �     �_�w� �     �    �  (�
  ��^  "  �    ����� v          �  X�  K�^  "  K    ����� 6          �  (�
  �_  "      ����� 6          �  S�  +�^  �  + !  �_�w�      �    �  �ǈ  +�_  	H  +  � �����           �� ��  �_�     @ ����           �� ��Ѐ �[� �P�     z��             �� zs�� �� �����    }\_      x O   �� >�.  �-�� .�   }���`     <     �x ?�~� �,��?  �  ����     >  >  �>7߁��� �,~7߂ ��  �?}�~      |  ������� �?���c��    ���     � �   ������ +������ (   ���     ��   ������� /��������,   ��     ��   � ���> /� �����~�h   ���     ���   �   ��� W� >��? P    ��� �8     ��   �   ?�  _�   �� @X    �  �0     >�    �   �  ���  7t @�    �  �p     p     �    �  ���  � @�       �`            ��   � �_��  � �@        �          @ ��  � �� �  � �`        �          @ `  � ����`  � ��  �     �          � p  � ����p  � ��  �     �         � ��  � ���@�  � ��  `                 ��  � �� L  � �  0                 ��  � �� 6  �                    ��  � o�� � � l                   ��� � _��� /� �       (           ���   ���@� _  ?�        p         0  �t>  ?�  w�>  ?`   � �   �         `  =����  ~�� ���  ~�   ��   �   ��    �  ����  ��  ���  �    p    �    @       ���� ���   w�� �     8         0       ��  ��x  �9�  � �       <            ��@  7��  p  4 @   �   �         0   ���  ���  �  |�    �  �     �   �   ��c��_��   c��`      �  �      `       ���?���    \?��     ?��              }������    ��       ���       ��     �������      ���        �         ?�      �������   @ �                          �������                                                                   Q Q  g�����0   �    �                         �������   @                           �����d   �     �                         n�������         D                        �������    �                         ��������  H �� 	      �                _�����`  � � �   ��              ��������  @ q���       8  @            ���  8���  ����    � p    �            ��0 �?��  > �  P   �  �              ���  ��  �        ��            /��  <'��  � 8<$     ��             [��   �3�� $ a� `��      ?               ��R  B 	���( �  � 9 
 @ ,  |        @     ���  � ���@�  � �  \  �        �     o�D  � ?� �D �  � �  � �       �     _��   ?� ��   � 8 �  �            ��H   ��� �   � @0 �  `            ��H   O��@H   H   0 �  0           �      ����    D   p �  8             �  `  !���$� t  "   p �               ��  �  �� l� ��    p s�             ��  ��  	�� X� ��� 	    p p        p     �     � �� ��� �  `p p              ��     �� �� �  �  @p                 �@H �L� ��@H 泀 �  �0 �� �     �@�  � �@@��� ��`D�3���  �8 �� �     ���  � �@� ����`D����B�  �8  a���      @� � �� ��� A_�� ��� Q`  >� ����    � � @@ ��� � ��#��� `  �����   � � @ ������ /� ���� 0  �������   �� �    �  ��� ����!��  �=���`      |    � ?�~`@���?� �y��  ��?�>`    >  >    � >�>����? ~�0�  ��ߟ `    <      � z@�/  ���z�b���  �^�_ `    x      � ��� W� ��P�X   z�� �     �    �  ��  W�   X   �����         �  ��� _�  X X   ����� �          �  s�  _�  � X   �_�w� �     �    �  (�
  ߀  " �   ����� 0          �  X�  ߀� "  �   ����� 0          �  (�
  [�� "  �   ����� 0          �  S�  [�  �  \ � �_�w� 0     �    �  �ǈ  [�@ 	H  \ � ����� 0          � ��  _��   X @ ���� 0          �� ��Ѐ _�� �P� X   z��  0           �` zs�� ��� ����� �  }\_  p    x O    �p >�.  ���� .� �  }���` p    <      �8 ?�~� ����?  � � ���� `    >  >   �߁��� ���7߂ �� � �?}�~ `     |   ��������/�߇��c��0  x��� �    � �    �������_�������@   ��� �    ��  @ �����������������`   �� �    ��  @ �@���>��`�����~��  � ����    ���  � �@  �����`>��?�  �  ��� ��     ��  � �`  ?� ��p  �� D�  �  �  ��     >�   � ��  � ��  7t E   @  �  ��     p    ��   � 	�� �  � I�  @     �            �X   � �� �  � ʀ                    ��  � ��� L  � �   0                 �  � ����&  � �                    �  � ����3  � �                    �� � W��@� � �        8           ��� � ��� 
� � �       p            ��@ � _�� @ � P   �    �         @  ��� � ��� � � �   �   �    �     �  ��X � ��X /� =@   �   �    @       ��$   2���@ � _  r�   x                 �� >  e��   S>  �     <��              =���� ���  �� �     ?   |     8      ��� '��  
� $    �   �             ���� 8���   �� 8�     �  �     �   �   �q��_�x  � q��` �    �  ?�      p      �������   ,�  @    ��             ��������   ��      ���       ��    ���������    ���        �         �      ���������     �                           }�������                                   �������                                    �������   @                             �������                                                                   Q Q  g�����0   �8  �                         �?���}�   @�  �                      ~�����d   �    @�                        n������       D                        ��������                            ���������  H@    	                        ^������`  �  �  B�  �     �             ���`���  B  �� !     �   @            ����/���   �0     � �� �            �������  1�� P      �               ��O���  ���    0 �            /��< <��  > <    � ��             [���  ���� $@�  ǐ     ? `              ��� B ����( 	� C� 
 @�  |  �      @     ���  � 7���A � � t A    �        �     m��  � �� � G  � 9 $�  8  �         �     _�   � � �  �� x �              ��  ?�  @ @ � � �            ��H   ��HH     � �  �           ��    /����    0  0 �  �            o�@ ` ����� t' �   0 �  `             ��  �
  ���� �*� �   p s�  p           ��  ��  K�� � ��� L  p p  8      p    ��     +�� � ��� h   p p             ��     7��@,� �  6   p                 ��H �L� ��@,H 泀    0 ��       �@�   �@��� ���XD�3�� @ 8 ��       ���   �� ��
���XD����J    8  a��       @�  � ��� M��0 ��� ]�  @>� ���     � � A  � #� � �� �#��� �  @����    � �   ������ � ����    @�������   �� �   �` ��� �� ` �!��  ��=����      |  � �@?�~`@��`?� �y��  ���?�?�    >  >  � �@>�>���`? ~�0�  ���ߟ �    <    � �@z@�/  ��`z�b���  ��^�_ �    x    � ����� _� ���P�`   z�� �     �   @ �� ��  ��  `   �����        @ �� ��� �� X `   ����� �         @ �� s�  �� � `   �_�w� �     �   @ �� (�
  ��� " �   ����� @         @ �  X� ��@ " � � ����� @         @ �  (�
 o�@ " p � ����� �         @ �@ S� o�@ � p � �_�w� �     �   @ �@ �ǈ �@ 	H ` � ����� �         @ �  �� �   ` � ���� �         @ �@ ��Ѐ_� P �P�` � z��  �          @ �` zs����h ������  � }\_ �    x O  � �p >�. ��t� .��  � }���`�    <    � �8 ?�~���9�?  ��  ������    >  > � �>߁����� >7߂ ���  ��?}�~�     | � ��������� ����c��   @x����    � �   �'������� �������  @ ���     ��   ���������3��������  @ ��     ��   ����>
���X�����~�     ���     ���   �  ������X>��? @   ��� �      ��   ��  ?� ��@,  �� U     �  �      >�    ��  � ��@.  7t V     �  �      p    ��   � /��   � l        �            ��   � ���   � �       8            ��  � ���	� � �        8            o�� � ����� � �        p             w�@ � ����` � �  �    `         @  ��  � ��@0 � @   �    �         @  ��� � ���  � � �   �   �    �     �  ��� � ߀ L � =�    p        @       ��� � 6���  6 � 7     8        0       ��� � i��� 	�/� �                   ��� ��}�@��_ � �       p            ��`> o��   > p     �� �         `   =���� 9���  �� ��      �  �      �  �   ��������  ��ƀ    p  ?       0      �����;���    o��:        �         8    {������x  � �� �    ���       ��    ���������   ���  @     �         �     ������{�  � �  �                        ���������                                   ���������                                }�������                                   �������                                   �������   @                            �������                                                                   Q Q  g�����0   �8  �                         �?���}�   @�  �                      ~�����d   �    @�                        n������       D                        ��������                            ���������  H@    	                        ^�������`  �      B�  �     �             ���������  B      !          @            ���������            �      �            ��������   �  P                       ��������  ��      �              /����?���   �0    ��               [���� ��� $@ ��      ?�               ���� A1���(  G�A� 
 @� 8 ~  �      @     ���� �����A � �<� A   ` �        �     m��` �?�� � x �0 $�  � � �        �     _���  ��� � �� �  � `             ���  o�� 	� �  @  �              ���   ���H   v     �             ��    ���� &         �              o�� ` ���� @ t' �    8 �               ��� �
  ��� � �*��    p s�              ��  �� _��  ���`   � p �      p    ��     ���  ����   � p �         �  ���    ��@� � p   p     �          @  ��H �L� ���@� 泀�   0 �� `      �@�    �@��� ����	��3��� @8 �� p      ���    �� �����D����T   8  a��       @�  � ��� S��� ��� T   >� ���     � � P  ��#� � �� #���    ����    � �   ������ �� ���    ������    �� �   �� �����  �!�   �=���       |   ��?�~`G�� ,?� �y�   ��?�<     >  >   ��>�>��� ,? ~�4   ��ߟ      <     ��z@�/ �� ,z�b��   �^�_      x     �����
�� X��P�     z��       �    �� �� 
�� X       ����          �� ��� 
�� X X      �����           �� s� �� X �      �_�w�      �    �� (�
 �� X "      �����           �� X� �� X "      �����           �� (�
 �� X "      �����           �� S� � X � �    �_�w�      �    �� �ǈ �� X 	H      �����           �� �� 
�� X       ����           �� ��Ѐ
�� X �P�     z��             �� zs���� , �����    }\_      x O   �� >�. �� (� .�    }���`     <     �� ?�~��� -�?  �   ����     >  >  ��߁����� 7߂ ��4   �?}�~      |  ��������+�� ���c��(   x���     � �   �������/�� �����,    ���     ��   �������S����������    ��8     ��   ����>_��������~�    ���0     ���   �  ���������? @  ��� �      ��   ��� ?� ?��@� �� 0     �  �      >�     ��� � O��@� 7t P     �  �      p  @  ��`  � �� ` � `   �   �          @  ��0  � ��� 0 � �   �   �          �  ��� � ���� � �    `        @       o�( � ��� � � �    p                w�� � 6���� V � 7    8               ��� � m���@ + � n                    ���� ����  ���       p            ���`�7�߀ 
`�8     �  �             ���������  ���     � �     �   �   ���FO�1?��� Gπq@     �0 �      @      ��y���}�@� ��΀ �    >  ?       8      ���?�1���    ~?�2       ��         0    =��������   ��       ���       ��    ��������   ��`      ?��        �     ��������     ?��                          {�������x  �      �                       ���������         @                       ������{�  �     �                        ���������                                   ���������                                }�������                                   �������                                   �������   @                            �������                                                                   Q Q  g�����0   �8  �                         �?���}�   @�  �                      ~�����d   �    @�                        n������       D                        ��������                            ���������  H@    	                        ^�������`  �      B�  �     �             ���������  B      !          @            ���������            �      �            ���������       P                       ���������                            /���������                              [��������� $@  �                         �����?����(  ��  
 @�  �   �            �����o����A  �p  A    �?�              m��������� �  8���  $�    �p         �     _��g����� �  ���  �  �              ������ �}�  @   �              ���0 ���H <@     ���            ��@  ����� p  �    �� @             o���d& ����� �t'�      �                ��� �* o��� ��*��      s�              ��� �� 7���   ���t     p        p     ���   ���  & ���2      p              ���    
���@ D �      8                 ��� �L�
���@ @ 泀
     8 ��       �@�   ��������� ��3��� @ x ��       ���   �� �����������    �  a��       @��  �@��� ����@��� �    �� ���     � � �  ���� � ��  ���� @   ����    � � @  ������� �� ��� `   ������    �� � @  ������_�� ��!�@   �=���       | @  ���?�~`/�� �?� �y�   ��?�`     >  >    ��>�>���� �? ~�   ��ߟ p     <      ��z@�/ ��� �z�b���   �^�_ p     x      �������� ���P��    z�� 0      �    �� �� W��   X    ����0          �� ��� _��  X X    �����0           �� s� _��  � X    �_�w�0      �    �� (�
 _��  " X    �����0           �� X� W��  " P    �����8           �� (�
 W��  " P    �����8           �� S� _��  � X    �_�w�0      �    �� �ǈ _��  	H X    �����0           �� �� W��   X    ����0           �� ��Ѐ��� ��P��    z�� 0            �� zs��� �������    }\_ p     x O    �� >�. ��� � .��   �}���``     <      ���?�~��� �?  ��   ����`     >  >   ���߁���_�� �߂ ��@   N?}�~�      |@  ���������� ���c��`   ����     � � @  ���������  �����@    ��� �     �� @  ����������������    ����     �� �  ����>��������~�    �����     ��� �  �� ������� ���=� @ @ ���       ��   ��X ?� ���@ � �� �      �        >�    ��� � 3���@ L 7t 3     0 �        p    ���  � 7���  & � 6                     ���  � o���  ; � l                   ���� ���� �� �        0            o��@�?���� @�0     �  �             w��0����� 0�`    � �         @   ���������@ ���      � �      �  �   �����r����   ��r�     x               �����Ǐ��߀  x��        |             �����w����   �t       ��         p    ����������  ��      ���        ��    ��������}�@� ���  �     ?�         �     ���������     �                           =���������                                 ���������                               ���������                                  {�������x  �      �                       ���������         @                       ������{�  �     �                        ���������                                   ���������                                }�������                                   �������                                   �������   @                            �������                                                                   Q Q  g�����0   �8  �                         �?���}�   @�  �                      ~�����d   �    @�                        n������       D                        ��������                            ���������  H@    	                        ^�������`  �      B�  �     �             ���������  B      !          @            ���������            �      �            ���������       P                       ���������                            /���������                              [��������� $@                             �����������(        
 @�       �            �����������A        A                     m�������� �   �   $�                      _������� �   p�  �   �                ���� o���   p   @   ���               ����������H  ��      �`              ���  g�����  �'�      �              o���`�����  o�'�       �               ����
����  ��*��      `s�              ��� �����  0���@     �p �       p     ���@ ����  `����     �p @             ���    _���@ @�P     �   �              ��� �L�����@ �泀�      ��P       �@�    �����G���� 	�3��  @  ��8       ���    ��� ������ ����       a�        @�   ���������  ���     � ��      � �   ���� � ���  #���     ���     � �    ����������  A���     ?�����     �� �   ������
���  P�!�
     /�=��        |   ���?�~e��  (?� �}�    G��?�      >  >   ��$>�>����  �? ~�    C��ߟ      <     ���z@�/��  �z�b��     A�^�_�     x     ������?��  ���P�@    @z���      �    ��@����� `�    ����        �  ��@������ `X�    �������         �  ��@s���� `��    ��_�w��      �  �  ��@(�
��� `"�    �������         �  ��@X���� `"�    �������         �  ��@(�
��� `"�    �������         �  ��@S���� `��    ��_�w��      �  �  ��@�ǈ��� `	H�    �������         �  ��@����� `�    ����         �  �����Ѕ?��  ��P�@    @z���            ���zs����  ������     @}\_�     x O   �� >�.%���  �> .��    @����c      <  !   ���?�~���  .?  ��    Q����      >  >   ���߁������  W߂ ��     .?}�~       |
   �����������  _��c��      ���      � �   ����������  /����     ���      ��   ����������� /�����     ��      ��   �����o���� ����l     ���      ���   �� ���s���� ��t  @  ���       ��   ����?� ����@ ��� �      � 0       >�    ���������@ �7t�      � `      p     ���  ����   �`     � �         @   ���� �����  ���     � �      �   �   ���������  ���      x        `      o��ӂ�������  S���       <              w���q������  <q�      � �             �����k����@  �l       ��         `    ����������   ��      ���        ��    ����O���߀   ���        ?�         �     �����������    �                           �����������                               ��������}�@�       �                       ���������                                  =���������                                 ���������                               ���������                                  {�������x  �      �                       ���������         @                       ������{�  �     �                        ���������                                   ���������                                }�������                                   �������                                   �������   @                            �������                                                                   Q Q    <�       � �       @                  �đ�      ;n        �                 >�>`      �� ��      @                  �����               @                ;��f     �l�      �                 L�?�_�     3��f      � @�               �������    @       �  �              g�����`    �   �     @                  ����?�   �   �`                        ;�����h   �    �                       �������                @              =�������                               [�������   $  ?�    @                  ��`?�v�  H��� �      �                n���o��@  � �p D�  @  �?�              }�������`  � ���  �  !  �p B       �     ��' p�� D ��� @   �              ����� @�}�     �             ��0 _�� <`  � ��� �           
��@  ���  p  � P �� @             ��` ��� 	 �t'�@   �               �� �
 k�� 
@��*��     s�              +�� �� 7��  3 ���t    @ p       p     ;�   �� �" ���2    p              W�    �� (�D �    8                  W�@ �L�� ( � 泀�@  8 ��       �@�    ��������	 ��3��  @ x ���      ���    ��� ����B�����  �  a��       @��  ��@��� ?߀P@���     �� ���     � �    ���� � _� R���� ` ������    � � @  {������ _������� @  ������    �� � @  _�������!�  �=���       |    [��?�~`/����?� �y0   ��?��     >  >    ��>�>��� �? ~�����ߟ p     <      ��z@�/ ��@�z�b��� �^�_ p     x      ��������H���P��    z�� 0      �    �� �� W��H  X    ����0          �� ��� _��  X X	 H �����0           �� s� _��H � X    �_�w�0      �    �� (�
 _��H " X    �����0           �� X� _��  " X	 H �����0           �� (�
 _��H " X    �����0           �� S� _��H � X    �_�w�0      �    �� �ǈ _��  	H X	 H �����0           �� �� _��H  X    ����0           �� ��Ѐ���H��P��    z�� 0            �� zs��@�������  }\_ p     x O    �� >�. �� �� .���� }���`p     <      [����~������  ��   ~���`     >  >   _��߁���O�߂ ��P N?}�~�      |@  {�������������c��`  8����     � � @  �������_� R �����` �� ����     �� @  ��������߀P������   ����     �� �  �����>���B����~�  �����     ��� �  ��� ������	 ���=� @ @ ���       ��   W�X ?� �� ( � ��  @    �        >�    W� � �� (�\ 7t      �        p    ;� � 7�� �& � 6                    +��  � o�� @ � l                   ���� ��� 
 �� �        0            ��@����  @��     �  `             �������  ���   @  @         @   �����x  ���� �    � �      �  �   ����r���   ��r�     x               ����ǎ���   X��       ? |             ����u���  ! 7�v B     ��         p    ��������  @ ��      ���        ��     ���������    ���        �         �      w�������   @ �                          /�������                                �������         @                         �������                                  �������                                   �������     @                             w�����@    �  �                          ~���      � @�                           /��o��      �                            �����       @                           �����      @                              ��o��       �                             ;���       @                                                          Q Q    <�       � �       @                  �đ�      ;n        �                 >�>`      �� ��      @                  �����               @                ;��f     �l�      �                 L�?�_�     3��f      � @�               �������    @       �  �              g�����`    �   �     @                  ����?�   �   �`                        ;�����h   �    �                       �������                @              =�������                               [�������   $        @                  ������v�  H�     �                        n������@  �  �  D�  @                   }��0��`  �  ��  �  !  �  B             ����o�� D �p @    ���         �     �������� @ ��     �`             ��ӂ ����  3��   � �  �           
��N  9��   �  y� P  0�              ���`��� 	 �t'�@   @�              ��`�
_�� 
@p�*�`     �s� �             +��������  �����    @ p `      p     ;�  ��� ������    p               W�    o�� (� � �                     W�� �L�'�� ( 3 泀d @   ��       �@�    ������3���	 "�3��  @  ��       ���    ���� �����B @����   <  a�        @�   �������߀P @���    >� ��      � �    ��C� ��� R ����  �� >���     � �   {������ ���� ���� �   _�����     �� �    _����� ��!�   O�=��       |   [�h?�~f���h?� �~@    ���?��     >  >    ��D>�>��� d? ~���� ���ߟ�     <   �  ��Bz@�/��@bz�b���  ��^�_�     x   �  ��A��󐂿��Ha��P��    �z���      �  �  �����_��H�`    �����        @  �������� �X`	 H ������         @  ���s���H��`    �_�w��      �  @  ���(�
��H�"`    ������         @  ���X�_�� �"@	 H ������         @  ���(�
_��H�"@    ������         @  ���S���H��`    �_�w��      �  @  ����ǈ�� �	H`	 H ������         @  �������H �@    �����         @  ��@��Ђ���H`�P��    �z���          �  ��@zs��@`������  �}\_�     x O �  ��@>�."��  a� .���� �}���a�     <   �  [�`?�~����� f?  ��    ������     >  >�  _��߁��� �߂ ��   N?}�~�      |	   {�?�������� ���c���   @���      � �   ��������� R _����  ��  ���      ��   ���������߀P _�����     ��      ��   ������u���B /�����   ���      ���   ��� ���%���	 ,��f  @  ���       ��   W�� ?� k�� (  �� h @   �        >�    W��� ��� (��7t �    � 8      p    ;�� ���� �
���      p             +��` �O�� @`�P    �  �         @   ������� 
 ���     � �      �   �   ��L�?��  L�9@      � �      @      ��3�����   ����    |        0      ������x  � ,���  �     |             ����g���   �h      ��         `    ���t���   t        ���        p     ���������  !  O�  B      ?�         �     ���������  @  �                           ���������                                   w�������   @                             /�������                                �������         @                         �������                                  �������                                   �������     @                             w�����@    �  �                          ~���      � @�                           /��o��      �                            �����       @                           �����      @                              ��o��       �                             ;���       @                                                          Q Q    <�       � �       @                  �đ�      ;n        �                 >�>`      �� ��      @                  �����               @                ;��f     �l�      �                 L�?�_�     3��f      � @�               �������    @       �  �              g�����`    �   �     @                  ����?�   �   �`                        ;�����h   �    �                       �������                @              =�������                               [�������   $        @                  ������v�  H�     �                        n�������@  �      D�  @                   }�������`  �       �  !      B             �������� D      @                      ���0��� @  ��      �               ��� _���   `   �  ���  �            
��������   ��  P  �`              ����&���� 	  3�'� @   �              ����
��� 
@ o�*�      s�              +��X����   �����    @  p       p     ;�  ?�� �8���@    �p�             W�@  �� (�`�    �   �              W����L���� ( �況� @   ��`       �@�    ������o���	 ��3��  @  ��0       ���    ���� �����B 	����     a�        @�   �������߀P ���    � ��      � �   ���� ��� R ���  �� ���      � �   {����������  ���    �����      �� �   _������ (�!�   �=��        |   [��?�~b���� X?� �s     '��?�      >  >   ���>�>���  \? ~� �� #��ߟ      <     ���z@�/��@ Zz�b��   !�^�_      x     ��ф�����H Y��P�      z��       �    �� ����H ��    @����           �� �����  �X�	 H @�����            ���s����H ���    @�_�w�       �    ���(�
���H �"�    @�����            ���X����  �"�	 H @�����            ���(�
���H �"�    @�����            ���S����H ���    @�_�w�       �    �� �ǈ��  �	H�	 H @�����            ��0����H ��    @����            ��P��Њ��H ؅P��     z��             ���zs����@ X�����    }\_      x O   ���>�.+��  Y� .� ��  }���f      <  "   [��?�~����� ^?  �     !����      >  >   _��߁���� +߂ ��   ?}�~       |   {����������� /��c��    ���      � �   ��������� R ����  �� ���      ��   ���������߀P �����    ��8     ��   ����������B �����   ���8     ���   ����������	 ����  @  ���p      ��    W��@?�W�� ( `��X @  �� �      >� @   W�0�o�� (�07tp   ���      p @   ;�� ���� ����    � �      �  �   +��� �2��� @��2�     x               ��S����� 
  ӆ��      <              ���q����   lq�       � �             ����k���   �l     ��         `    ������x  � ��  �    ���        ��    ���������   ���       ?�         �     ���������    ?�                           ���������  !      B                        ���������  @                               ���������                                   w�������   @                             /�������                                �������         @                         �������                                  �������                                   �������     @                             w�����@    �  �                          ~���      � @�                           /��o��      �                            �����       @                           �����      @                              ��o��       �                             ;���       @                                                          Q Q    <�       � �       @                  �đ�      ;n        �                 >�>`      �� ��      @                  �����               @                ;��f     �l�      �                 L�?�_�     3��f      � @�               �������    @       �  �              g�����`    �   �     @                  ����?�   �   �`                        ;�����h   �    �                       �������                @              =�������                               [�������   $        @                  ������v�  H�     �                        n�������@  �      D�  @                   }�������`  �       �  !      B             �������� D      @                      ��������� @                            ��������   �    �       �            
��������    p   P   �               ��������� 	  ��� @                     ����
/��� 
@ �:�      s�@              +��������   ���     @ pp       p     ;�� u��� � 3���     p              W��  ��� (� F�9     8                 W���L��� (  �泜� @   p��        �@�    ������?���	 �3�@  @  ����       ���    ���!� ß���B !��ߠ    �  `�        @�   ���G���_�߀P G���@    �� ��      � �@   ���O� �?�� R O���0  �� ����      � �    {�����/���� ��     �����      � �    _������ �!�   �=��        |   [��?�~���� ?� �     ��?�      >  >   ���>�>���  ? ~� �� ��ߟ8      <     ���z@�//��@ z�b��   	�^�_      x     ���������H ��P�     z��       �    �����7���H 4     ����           ���������  ,X 	 H �����            ���s����H ,�     �_�w�       �    ���(�
���H ,"     �����            ���X����  ," 	 H �����            ���(�
���H ,"     �����            ���S����H ,�     �_�w�       �    ����ǈ���  ,	H6 	 H �����            ��������H ,6     ����            ����Ы���H �P�     z��             ���zs����@ �����   }\_      x O   ���>�.K��  � .� �� }���8      <     [��?�~����� 
?  �     ����8      >  >   _��߁���� ߂ ��   ?}�~0        |   {����������� ��c��    ���p      � �    ��������� R ����  �� ���`      ��    ���G���_�߀P ���@    ����      ��@   ���!��Ɵ���B 5��Ơ    �����      ����   �����������	 ����  @  �����      ����   W��H?��� (  ̾�� @   p�       @>�    W���&��� (� w7tg     8�       0p    ;�Ɂ����� � )���      <             +���s�3��� @ {�4      � �         0    ��������� 
  ���       ��       � �    ���p?���   p@        ���        p     ���������    O�       ?�         �     �������x  �  �   �                       ���������                                ���������                                 ���������  !      B                        ���������  @                               ���������                                   w�������   @                             /�������                                �������         @                         �������                                  �������                                   �������     @                             w�����@    �  �                          ~���      � @�                           /��o��      �                            �����       @                           �����      @                              ��o��       �                             ;���       @                                                          