��`  |J� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         ����������������������������������������������������������������������������������������������������������������������������������������������������������������������� �                                       ������������������������������������������������������������������������������������������������������������������������������ ����������������������������������������������������������������������������������������������������������������������������������������������������������������������� �������������������������������������������                                       o���������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������    �       �                      p �������������?���������������������������������������������������������������������������������?�����������������������������   �       � � �                  p �������������?�������������������������������������������������������������������������������?���������������������������   `      �   0     0             p ���������������������������������������������������������������������������������������������������������������������������   `          `     `             p ������������������������������������������������������������������������ ���������������������������������������������������   0@      �   �     �     @      p �����Ͽ��������������������������������������������������������������� �������������Ͽ����������������������������������   `       �  ��     �    @      p ������������������ �����?����������������������������������������������  �������������������������� �����?�����������������   � �� � ?��� ��    @�     p �����?�>�y���}��������??���������������������������������������������  ������������?�>�y���}��������??����������������  ��ǁ�� ����?��   �@�     p �����?�8~9���<��~���>������?�������������������������������������  �������������?�8~9���<��~���>����������������  ����~ ������a�   �@��    p ������� �?���9��>�����������������������������������������������    ������������� �?���9��>�������������������   �o���=� 8�7c��     �     p ��������D�~��q��|��<Ȝ|<���������������������������������������������    ?��������������D�~��q��|��<Ȝ|<�����������������   �o��8q� 1�>��     �     p ��������	��s��sǎ|��|�<�|���������������������������������������������    ?��������������	��s��sǎ|��|�<�|�����������������   �8�0� 3�|Ä    8 �     p ������������������|�<{����������������������������������������������    ������������������������|�<{������������������   3�q�80c<1�cy��    8�     p ��������3�#��Ϝ��8����~����������������������������������������������    ��������������3�#��Ϝ��8����~������������������  �7�a�81�xc�<c�>    p�     p ������g�s������x�Ü������������������������������������������������    ������������g�s������x�Ü��������������������  0w�8pg�xg����    p �     p ������ψ�GǏ�y����9�|8��������?��������������������������������������    ������������ψ�GǏ�y����9�|8��������?����������  0fð0�n������     p�'      p ������ϙ�<O�����?9�<�<��������??�������������������������������������    ������������ϙ�<O�����?9�<�<��������??���������  0�9�pa�|��<���     � �"      p �������1�8����O3��~y�8���������>��������������������������������������    �������������1�8����O3��~y�8����������>����������  3�1�`g`�0���y�8    �A      p �������3�p�����3��y�y�����������������������������������������������    �������������3�p�����3��y�y��������������������  �?�0��~`�a���0<    �@�     p ������c� ���p3���y�����������������������������������������������   p������������c� ���p3���y��������������������  �`�@<�@a����   �A      p ��������	��?���xg���>�������?���������������������������������������   ���������������	��?���xg���>�������������������                    �    ��      p ������������������������?�����?����������������������������������������   �������������������������������?������������������                         � ��      p ������������������������������?����������������������������������������   ��������������������������������������������������                         � ��      p �����������������������������������������������������������������������   p��������������������������������������������������                         � C      p �����������������������������������������������������������������������    ��������������������������������������������������      8                   � A      p �����������������������������������������������������������������������    ��������������������������������������������������      p                     "      p �����������������������������������������������������������������������     ��������������������������������������������������      �                     "      p ����������������������������������������������������������������������      �������������������������������������������������      �                     "      p ���������?�������������������������������������������������������������      ���������������?����������������������������������                                  p �����������������������������������������������������������������������     ��������������������������������������������������   � �   0`   � `               p �����<�����ϟ����?���������������������������<�����ϟ����?�����������     ����������<�����ϟ����?�������������������������   � �   0   � `        
      p �����<�����������?���������������������������<�����������?�����������    ����������<�����������?�������������������������   f �   0   � `        
 �    p �����������������?��������������������������������������?�����������   �����������������������?�������������������������   <<�3<�>g��>��|x�       @�    p �������3���p��fa����������������������������3���p��fa�����������   �?������������3���p��fa�������������������������   f�3f ٻlٳf�fͶ       @�    p ������3̙�&D�&L��g�2I�����������������������3̙�&D�&L��g�2I�������   �?�����������3̙�&D�&L��g�2I���������������������   f�~�3o�?f��f��      8 ��    p ������3��'̐0���2�9������������?�����������3��'̐0���2�9�������   �?�����������3��'̐0���2�9���������������������   f�`�3l0f̀f�f      8 ��    p ������3��'̓�ϙ�2�?������������?�����������3��'̓�ϙ�2�?��������  ������������3��'̓�ϙ�2�?����������������������   f�fٳl�3f͘fͶ      8 ��    p ������#��&L�9̙�2g�2I�����������?�����������#��&L�9̙�2g�2I�������   ������������#��&L�9̙�2g�2I���������������������   <|<�3g�>��|x�      p ��    p ������Ã���0̘y���3������������?������������Ã���0̘y���3���������   ������������Ã���0̘y���3�����������������������                           p  �    p ���������������������������������������������������������������������   �������������������������������������������������                           p  �    p ����������������������������������������������������������������������   ��������������������������������������������������                           �� ��    p ���������������������������������������������������������������������   ��������������������������������������������������                           �  �    p ���������������������������������������������������������������������   ��������������������������������������������������                           � ��    p ��������������������������������������������������������������������  ��������������������������������������������������          0  ��    0      � � �    p ���������������>������������?������������������������>�������������   ���������������������>���������������������������         `` �     0      � � �    p ���������������?�������������?���?���������������������?��������������   ���������������������?����������������������������         `` �     0      �   �    p ���������������?�������������?������������������������?��������������?   ���������������������?���������������������������   q��x�ps����?�0      �   |    p ������1��a��1�c�0�p�������������������������1��a��1�c�0�p���������?   ������������1��a��1�c�0�p�����������������������   �6l��`fl���ٰ      �   |   p �����$ɓ3�L����I�>I&O�����������������������$ɓ3�L����I�>I&O��������?   �����������$ɓ3�L����I�>I&O���������������������   cl��`fl͘϶߰      �   |   p ���������@����2g�0I O���������������������������@����2g�0I O�������    ���������������@����2g�0I O����������������������   3l��`fl͌ٶ�0      @   >   p ��������?�O����2s�&I'���������������������������?�O����2s�&I'��������    ��������������?�O����2s�&I'����������������������   �6l�3`flͶٶـ      �   >    p �����$ɓ3�̟���2I�&I&�����������������������$ɓ3�̟���2I�&I&��������   �����������$ɓ3�̟���2I�&I&����������������������   q��x0c�͜϶�0      �   >    p ������3���Ϝ3�2c�0I0�������������������������3���Ϝ3�2c�0I0����������   �?�����������3���Ϝ3�2c�0I0�����������������������               �         �   �   p ������������������?��������������������������������������?������������   �������������������������?�������������������������              �         � � �   p ��������������������������������������������������������������������   ��������������������������������������������������                          � @     p ����������������������������������������������������������������������   ��������������������������������������������������                           p         p ���������������������������������?��������������������������������������   ����������������������������������������?����������                             @      p ������������������������������������������������������������������������   ���������������������������������������������������                             ��      p ����������������������������������������������������������������������� ����������������������������������������������������                            ����     p �������������������������������   ��������������������������������������������������������������������������������������������                            ����     p �������������������������������   ��������������������������������������������������������������������������������������������                            � ��     p �������������������������������� ��������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������   ��                     0           p ����������������������������������������������?�������������������������������������������������������������������������������   ��     �         0     0           p ����������������������������������������������9?�����?�������������������������������������������������������������������������   ��     �         0     0           p ����������������������������������������������9?�����?�������������������������������������������������������������������������   ��8�|��f�����9�sǏ9�6y��Ǐ9�   p ����������������������������������������������90���c�a���8p�Ɇd~8p��������������������������������������������������   �كm�3v���f��m�30flٳ06͛lٳ0   p ����������������������������������������������&|�g̉3'�L�?�g�ϙ�&L��2d��&L��������������������������������������������������   �ߟ1�?f���f���m�30g��06͛���   p ����������������������������������������������? `���0'�L�?3��Ϙ�L��2d�s�L�������������������������������������������������   ��3�0f��f�͛m�30f�06͛ ��    p ����������������������������������������������?'��ϙ3��L�?2d��ϙ��L��2d�3�L��������������������������������������������������   �ٳm�3f��3n�͛m�30flٳ0ͻlٳ0   p ����������������������������������������������?&L�g̙3'�̑?2d�g�ϙ�&L��2D��&L��������������������������������������������������   ��8�fg�>���l��cǏ1�x�Ǐ1�   p ����������������������������������������������?0��ᙘg���?3���8p���8p��������������������������������������������������                                    p �������������������������������������������������������������������������������������������������������������������������������                          p          p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������    ?�����������������������������    p �������                            �������������������������������������������������������������������������������������������    ?�����������������������������    p ������������������������������������������������������������������������������������������������������������������������������    ?�����������������������������    p ������������������������������������������������                           ��������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    ?�����������������������������    p �������                           �������������������������������������������������������������������������������������������    ?�����������������������������    p ������������������������������������������������������������������������������������������������������������������������������    ?�����������������������������    p ������������������������������������������������                            ��������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������              �o߿   ` 6          p ������������������������������������������������������������� @���������������������������������������������������������������             c1�  ` 0 �        p ���������������������������������������������������������������|�������������������������������������������������������������             c1�  ` 0 �        p ���������������������������������������������������������������|�������������������������������������������������������������        3�9�c1���6��        p ������������������������������������������������������c��q����|a�p�������������������������������������������������������        6��6��c?3lٶ홀        p ������������������������������������������������������'�L�$�0�������&If������������������������������������������������������        3���1�3o�6���        p ��������������������������������������������������������L�����|���'�2������������������������������������������������������        �1����1�3l6́�        p ����������������������������������������������������$�g�L�y����|�����2~������������������������������������������������������        �v��6��1�3lٶ͙�        p ����������������������������������������������������$�'�L�$����|���&I2f������������������������������������������������������        q�1��c����6��        p ����������������������������������������������������s��q���N~a�p�3������������������������������������������������������                          �        p ������������������������������������������������������������������������������������������������������������������������������                                   p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p ���������������������������������������������������������������������������������������������������������������������������������������������������������������������� ��                                      ?����������������������������������������������������������������������������������������������������������������������������� ����������������������������������������������������������������������������������������������������������������������������������������������������������������������� �������������������������������������������                                       ��������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         ������������������������������������������������������������������������������������������������������������������������������