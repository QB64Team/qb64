�bt  @  ���>��00��>  ��@@��  ����  ���  �    ���   �� � ���G��6��?������?�������>��  �����        ���>��00��>"�"����EDED����ğ��"�2������  @��   �� � ���G��6��?������?�������>��  �����        ���>��00��>  ��AED���FG�Gď������������PP���
��#����h.�<���2r���8<|x���>�?�������>��  �����        ���>��00����  ����@@����@@�������������������� ����� ����@ ���� @����  ���� 0 ����� ����        ��    �������?�?��  ��   �F��  ���  ���  ���  PP�  ���   0�    �    �N� ����  ��  ��  �        ��    �������?�?��  ��  �����  @�B��  ���   0�    �    @�                    ��  �����  ��  ��  �        ��    �������?�?��  ��    ���   ���    @�                                            ��  �����  ��  ��  �        ��    �������?�?��  ��    ��    ��                                                    ��  �����  ��  ��  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      