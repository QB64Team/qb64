�i  $(� k 8                       8                       ?                       8                       G                       G                       |�                      D                       ��                      ��                      ��                     �                       ���                     ���                     ��>                     ��                      ���                     ���                     ���                    ��                     G���                    D���                     >                    D >                     ?���                    ?��                    8���                   8 �                    ~����                  z�?��                   $�                                         >���                   <���                   R >�                    �                   ? ?���                  = >��                   �p                                        ����                  ����                  )  �                     �                  � ��                  � �                  	  �q�                     p                  � ���                 @ ���                 �  8                                       �  ��                 @  �                 �  ��                     �                 �  ��                 �  ��                 
@   p9�                     8                 �   ��                �   q��                
@   0                                      �   ��                �   ?�                    ��                     �                �   ��                �   ��                     83�                     0                �    ?��               �    9��               �    `                �                     �    ��               �    ?�               �    Ø                �     �                �    ��                �    ��               H     0f                @      `                �     ?�                �     3�               H     �               @                      ~     ��               z     �               �     �`                                      ~     ��               z     ��               �      a�                      �               ?      �               =      g�               R      f                      `               ?      �               =      �               R      �                                    �     ��              �     �              )      �`                                    �     ��              �     ��              )       a�                     �              �      �              @      g�              �      f                      `              �      �              @      �              �      �                                   �      ��             �      �             
@      �`                                   �      ��             �      ��             
@       a�                     �             �       �             �       g�                     f                      `             �       �             �       �                     �                                  �       ��            �       �            �       �`             �                     �       ��            �       ��            �        a�             �        �             �        �             �        g�            H        f             @         `             �        �             �        �            H        �            @                      ~        ��            z        �            �        �`                                   ~        ��            z        ��            �         a�                      �            ?         �            =         g�            R         f                      `            ?         �            =         �            R         �                                 �        ��           �        �           )         �`                                 �        ��           �        ��           )          a�                     �           �         �           @         g�           �         f                      `           �         �   �       @         �   �       �         �  p                     p       �         �����       �         ����       
@         ����                  ���       �         �� �       �         �� �       
@          a����                  � �       �          � �       �          g�                   ���                   @         �          � �       �          �                   ?���                             �          � �       �                   �           ����        �                     �           � �       �           � �       �           ?��t        �                      �           ��r        �           ��r�      H           ( �        @                      �           � ��       �           � ��      H           )  w        @                     ~           � v        z           � 7        �           )                                ~           � 9�       z           � ?�       �           )  p                      0        ?           � A�       =           � ߠ       R           )   @                             ?           � `       =           � `       R           )  	�                    @       �          � �       �          � �       )           )                               �          � `       �          � �       )           )                               �          � `       @          � 7�       �          )                                �          � �       @          � �       �          )  p                           �          � `       �          � p       
@          )  �                            �          � �       �          � �       
@          )                               �          �        �          � �                  )                                �          �  �       �          � �                  )   �                     �       �          � �       �          �  �       �          )   `        �             @       �          �  �       �          �  �       �          )  �        �             �        �          �         �          � ~�      H          )           @                      �          �  9�       �          �  y�      H          )   '        @             !        ~          �  t        z          �  7�       �          )                                 ~          �  0        z          �  ?        �          )   p                      0        ?          �   �       =          �  ��       R          )   @                              ?          �  �       =          �  o�       R          )                                �         �  @       �         �  �       )          )                                �         �  @       �         �  �       )          )                                �         �  �       @         �  �       �         )                                �         �  �       @         �  �       �         )                                �         �  �       �         �  �       
@         )   �                    �       �         �  �       �         �  �       
@         )   �                     �       �         �  �       �         �  �                 )    �                     �       �         �  |       �         �  D                 )    �                     D       �         �   �       �         �  �       �         )    �        �             �       �         �   �      �         �   �      �         )    ��      �             �       �         �   � ��     �         �   � ��    H         )    ��      @             �        �         �   {       �         �   C       H         )    ����     @             @        ~         �    >      z         �          �         )    ���                          ~         �   �>      z         �   �      �         )   ����                   �      ?          �  ��>      =          �  �       R         ?  �����                  �       ?            ���      =            �        R         ?�������                 �         �         ������     �         � �       )         q����� ��                �          �        ����       �        � �       )         �����                   �           �        ?����         @        .� �         �        ���                                �        ?���          `        .��          �        ��                                 �       ?��           �        .��           
@       �p                                   �                   �                            ��                                   ��  � �             ��  �              ���������             �                     �������             ������               �����������             ?������               ����������               �  �  �              ���������               �  �                 �������                      �              ��������`                                      ��������               ������                �  �                                         �  �                  �  �                                                                 �                                              �                                              �    0                 �����                 �                                             ������                                        ������                                         �    <                                        �    4                                                                                                                                