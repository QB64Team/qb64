�,b  ��Q Q  g�����0   �    �                         �������   @ ?�                        ����d   ��� �      ?�                 n��  ��       D    ���                �������   c��      ?�              ���<���  H����	     `�               _�p(/�`  �~(0�  �� �             ��� @���  @�H�    � 0 @            �� @ q��  g�
H �    � �  �           �\ @ ��  � @ = P     �              �� p �� � p �   @ �             /�` p ?� p p   � �  �            [�� p �� $� p �    �               ��  p  ���(	� p �
 @  �  0           ��  p  w��@  p  �   �             o�  p  ;� �&  p  x�   �             _�  p  7� �l  p  6�   �             ��  p  �� X  p   @   �             ��  p  ��@�  p  �  @  �             ~   p  ?��0  p  @  �  �  �           @  gv  ���`  ww  �  �  �  �         � ��  �z  ��  �z�      s�   �     #"     ��  ��  ��  ��� `    p   �     p   @ �       ���  ��� �    p   `           �        ���  �   �         `            �   �L�  W�   泀  �    ��  0     �@�   �  ���  _�  �3�  X    ��  0     ���   �  � �  k�  ���  l     `        @   �  ���  +�  ���  l   � �      � �   �  � �  /�  ���  ,   ��      � �   �  ���  �  ��  6   ���      � �   �  ���  �,  �!�  6   ?=�~        |   �  ?�~  �,  ?� �     >�>      >  >   �  >�>  �,  ? ~     |�ߟ      <     �  z@�/  �\  z�b�      }^�_      x     �  ��� 
�X  ��P�     z��       �    �  ��  �X        ����          �  ���  �X  X      �����           �  s�  �X  �      �_�w�      �    �  (�
  �X  "      �����           �  X�  �X  "      �����           �  (�
  �X  "      �����           �  S�  �X  �      �_�w�      �    �  �ǈ  �X  	H      �����           �  ��  �X        ����           �  ��Ѐ �X  �P�     z��             � zs��  � z���      �\_      x O   � ��.@ �, � .@   ���߀    �     � ��� �, �  �   �����    �  ?�  � __���� �, __� ��   ?�}��      |�  �}/���= �}��c��   ����~    |� �<  ������@+������@( �����  ���  ��������/��������, ���� ���� �_O�������_������� ������  ��� � ��> ���><w�	�� ���p �  ��� � �  �� <p ��� ?� ��� �� >� �� �  �  �  �  >�  � ��� � ���� t �� �  �  �  �  p  � �π     ��� ��    �� �      �  �      � ��      ?߀�      � �      �  �      � �X      �� |      ?� �      �         � 0      ���8      �  �      �         � 0      ���0      �  �      �         � ��      ��@�      �  `                  ��      �� L        0                  ��      �� 6                          ��      o��       l                    ��      _���     �        (           ���     ���@�    �        p         0  �`    �  `    `   �     �         `  =��    �� �    �   �    �   �     �  ��    	�  �    	    p    �    @       ��    7��   v    7     8         0       ��   ��x  �9�   � �       <            ��`  7��  p  4 @   �   �         0   ���  ���  �  �    �  �     �   �   ��c��_��   c��`      �  �      `       ���?���    \?��     ?��              }������    ��       ���       ��     �������      ���        �         ?�      �������   @ �                          �������                                                                   Q Q  g�����0   �    �                         �������   @                           �����d   �     �                         n�������         D                        ���� ���    �                         ��������  H �� 	      �                _��  ��`  �    �   ���              ���� ����  @ s� �     �  @            ����G����  ��G��    � p�  �            ��~
H??��  ~
H?  P   �� �             ���@���  �@�     �              /��p ���  �p�    �              [�� p ;�� $ o p z     �              ��� p ��( \ p �
 @   �             ��� p ���@� p �  @ �             o�` p _� �p p `�  � �  �            _�� p �� �� p ��   �  @            ��� p ��� � p � @  �               ��  p  ���@  p  �     �             �  gv  u���  ww  v     �              �  �~  3���.  �� 2     �              ��  ��  �� ,  ���      p              ��  ��  �� X  ���       p        p     �0     	�� �  ��� 	�  @  p              ��  � � �� �  ��� �  @  � �       � �    �` �L� ��p �� �  �  ��       �@�    �@ ��� �` �3� @  �  �� �     ���    �@ � � _�` ��� `  �   ` �      @    �� ��� ?�� ���     � �  �    � �    �� � � ?�� ���     ��  �    � �    �� ��� �� ��    ���  �    � �    �� ��� ��� �!� �   ?=�~  `      |    �  ?�~  ��� ?� �  �   >�>  `    >  >    �  >�>  ��� ? ~  �   |�ߟ  p    <      �  z@�/  ��� z�b�  �   }^�_  p    x      �  ��� ׀  ��P� �   z��  0     �    �  ��  _�    X   ���� 0         �  ���  _�  X  X   ����� 0          �  s�  W�  �  P   �_�w� 8     �    �  (�
  W�  "  P   ����� 8          �  X�  W�  "  P   ����� 8          �  (�
  W�  "  P   ����� 8          �  S�  W�  �  P   �_�w� 8     �    �  �ǈ  _�  	H  X   ����� 0          �  ��  ߀    �   ���� 0          �  ��Ѐ ׀  �P� �   z��  0           � zs��  ���z���  �   �\_  `    x O    � ��.@ ���� .@ �  ���߀ `   �      � ��� ����  � �  ����� `   �  ?�   ��__�������__� ���  ?�}�� `     |�   ��}/���=/��}��c��0  ����~ �   |� �<   �E�����C�E�����C` �������  ��� @ ����������������` ������  ����@ �O������߀������� �������   ��� �� �>���>>�������  �  ��� �    �� >� �|� ?� ���� >� ��  �  �  �    >�  � �9� � ῀?� t ��  �  �  �     p  � ���     ��� ��    �  @                  ��      w� _      w�                     ��      w�� n      w                     �      n���.      o                     �      O���      L         8           ��      ���@      �         8           ���     ��� �     �        p            ��@    O�� @    P   �     �         @  ���    ���  �    �   �    �    �     �  ��P    	?��X    	@   �    �    @       ���    ���@ $        x                 ��    d��   S    e     <                =���  ���  �  �         |            ��0  /��  
0  (    �   �             ���  8���   �  8�     �  �     �   �   ���ǿ�x  ����� �    ~  ?       p      �������   l�  @    ��             ��������   ��      ���       ��    ���������    ���        �         �      ���������     �                           }�������                                   �������                                    �������   @                             �������                                                                   Q Q  g�����0   �8  �                         �?���}�   @�  �                      ~�����d   �    @�                        n������       D                        ��������                            ���������  H@    	                        ^������`  �  �  B�  �     �             ���`?���  B �� !     �   @            ���  7���     8     � ��� �            ��������  1�� P    ?�8               ��O$y��  ��'��    0�             /��8H��  >H>@   ���              [���@��� $@�
H�    � `             ����@ ����( �@� 
 @� �  �           ��� p 7���A  p t A   �             m�� p �� � N p 9 $�  0 �              _�8 p � � � p �� @ �              ��` p ?�p p @ @ � �  �            ��� p ���H � p �    �  @           �� p ����� p �    �  @           o�� gv  ����� ww  �     �               ��  �z  ���� �z� �     s�        #"     ��  ��  [��   ��� \    p  (      p    ��     +��   ��� (     p             ��  �   5��@,  ��� 6                     ��  �L� ��@,  泀      ��       �@�   � ��� ���X �3�  @   ��       ���   � � � 
���X ��� 
       `        @   � ��� ���0 ���    @ � �      � �   �  � � � � ��� �  @ ��      � �   �� ��� � � ��    @ ��� �    � �   �` ��� �� ` �!� �  � ?=�~ �      |  � �@ ?�~ �� ` ?� � �  � >�> �    >  >  � �@ >�> ��` ? ~ �  � |�ߟ �    <    � �@ z@�/ ��` z�b� �  � }^�_ �    x    � �� ���� � ��P�@   z��  �     �   @ �� �� _��  `   ���� �        @ �� ��� �� X `   ����� �         @ �� s� �� � `   �_�w� �     �   @ �� (�
 _�� " @   ����� �         @ �� X� _�� " @   ����� �         @ �� (�
 �� " `   ����� �         @ �� S� �� � `   �_�w� �     �   @ �� �ǈ �� 	H `   ����� �         @ �� �� � �  @   ���� �         @ �� ��Ѐ� � �P�@   z��  �          @ �@zs�� ��`z��� �  � �\_ �    x O  � �@��.@�� `� .@�  ����߀�   �    � �@����� `�  ��  �������   �  ?� � �`__������ `__� ���  �?�}���     |� � ��}/���=�� �}��c���  `����~    |� �<  �������E�� �����e�  {�����   ���  ������������������   ����   ����  �O���������G������   ?�����    ��� �  � ���>{���� ��z @>  ��� �     �� r  ��� ?� ���@'� >� �     �  l      >�  d  ��� � ���@� t �     �  ,      p  $  ���    ��� �    �                     ��     ��� �    �        8            ���     ����    �         p            o��    �����    �         `            w�`    ���`    `  �     �         @  ��0    ��@0    @   �    �         @  ���    ���  �    �   �    �    �     �  ���    �߀ L         p         @       ���    '���  2    &     <         0       ����   O��� �   L        8            ���  ��}�@��  � �       p            ��8  ��   8  `     �  �         `   =���  y���  �  y�      �  �      �  �   ��������   q��     >  >       0      ����?���    �<       ��         8    {������x  � �� �    ���       ��    ���������    �   @     �         �     ������{�  � �  �                        ���������                                   ���������                                }�������                                   �������                                   �������   @                            �������                                                                   Q Q  g�����0   �8  �                         �?���}�   @�  �                      ~�����d   �    @�                        n������       D                        ��������                            ���������  H@    	                        ^�������`  �      B�  �     �             ���������  B      !          @            ���������            �      �            ���������   �  P                       ��������  ��      ?�              /���  ?���     0    ���               [�������� $@ ��     �0               ����@1���(  G�C� 
 @� 8�  �           ����@����A �@<� A   `�             m��pp?�� � xp0 $�  �� �             _���p ��� � �p� �  � p             ��� p g�� �p �  @  �              ��� p ���H  p r     �             �� p 	���� . p 9     �             o�� gv ���� X ww �      �              ��� �z  �� � �z�@    @ s� �      #"     ��` �� _�� p ���`   � p �      p     ��@    ?�� ` ���    � p �            ���    ��@� � p         �          @  ��� �L� ���@� 泀�     �� `      �@�    � ��� ����	��3� � @  �� p      ���    � � � S��� ��� T      ` 8       @   � ��� S��� ��� T    � � 8     � �   �� � � /��  ��� ,    ��      � �   �� ��� +��  �� (    ���      � �   �� ��� ��  �!� 6    ?=�~        |   �� ?�~ �� , ?� �     >�>      >  >   �� >�> �� , ? ~     |�ߟ      <     �� z@�/ �� , z�b�     }^�_      x     �� ���
�� X ��P�     z��       �    �� �� 
�� X       ����          �� ��� 
�� X X      �����           �� s� �� X �      �_�w�      �    �� (�
 �� X "      �����           �� X� �� X "      �����           �� (�
 �� X "      �����           �� S� � X � �    �_�w�      �    �� �ǈ �� X 	H      �����           �� �� 
�� X       ����           �� ��Ѐ
�� X �P�     z��             ��zs�� �� ,z���     �\_      x O   ����.@�� ,� .@   ���߀    �     ������� ,�  �   �����    �  ?�  ��__������ __� ��4   ?�}��      |�  ��}/���=�� }��c���   ����~   |� �<  ��������� �����   �����   ���  ������������������   ����   ����  �G���������������   �����     ����  � ���=����� ��}� @  ����      ���  ��x ?� ���@� >� �     � �      >�  �  ��� � ���@� t �     � �      p  �  ��`    ��� p    �   �    �          �  ��     ��� 0    �   �    �         �  ���    ����    �    @         @       o�(    ��� �    �    p                 w��    6���� V    7    8                ���    m���@ +    n                     ���   ����  �  �        p            ���`  7�߀ 
p  8     �   �             ����  ����  �  �     �  �     �   �   ���F  1?��� G� �@     �  �      @      ��y���}�@� ��΀ �    >  ?       8      ����1���    ~�2       ��         0    =��������   ��       ���       ��    ��������   ��`      ?��        �     ��������     ?��                          {�������x  �      �                       ���������         @                       ������{�  �     �                        ���������                                   ���������                                }�������                                   �������                                   �������   @                            �������                                                                   Q Q  g�����0   �8  �                         �?���}�   @�  �                      ~�����d   �    @�                        n������       D                        ��������                            ���������  H@    	                        ^�������`  �      B�  �     �             ���������  B      !          @            ���������            �      �            ���������       P                       ���������                            /���������                              [��������� $@  �                         �����?����(  ��  
 @�  �   �            ����,o����A  ,p  A    �Ӏ              m����G���� �  8�O�  $�   �p               _��g�@���� �  ��O�  �  �              ����@�� �@}�  @   �              ���0p���H <p@     ���            ��@p����� pp�    �� @            o���gv ����� �ww�      �               ��� �z o��� ��z��      s�        #"     ��� �� ���   ���T    
 p (       p     ���   3���  . ���2      p              ���    ���@ L �      0                 ��� �L�
���@ X 泀
       ��       �@�   ��������� ��3�� @ @ ��       ���   �@� �����P����    �  `�       @ �  �@�������`����    �� ��     � � �  ���� ���  ����@    �� �     � � @  �������� ���`    ��� �     � � @  ������_�� ��!�@    ?=�~ �       | @  ���?�~ ��� �?� � �    >�> `     >  >    �� >�> ��� �? ~ �    |�ߟ p     <      �� z@�/ ��� �z�b� �    }^�_ p     x      �� ������ ���P��    z�� 0      �    �� �� W��   X    ����0          �� ��� _��  X X    �����0           �� s� _��  � X    �_�w�0      �    �� (�
 _��  " X    �����0           �� X� W��  " P    �����8           �� (�
 W��  " P    �����8           �� S� _��  � X    �_�w�0      �    �� �ǈ _��  	H X    �����0           �� �� W��   X    ����0           �� ��Ѐ��� ��P��    z�� 0            ��zs�� ��� �z��� �    �\_ p     x O    �����.@��� ž .@�   ���߀`    �      �����ѿ�� ��  ۠   o�����`    �  ?�   ���_����_�� �_� ��@   ?�}���    ?  |�@  ���/���?�� ���c��`   >���~�    <� �>@  ���w�����  �����@   8���>�    0��@  �S���������������    ����     ���  �g���������������    ����	�     ����  �� ���}���� � ���� @ @ ���       ��	   ��\ ?� :���@ � >� z�      �        >�    ��� � 3���@ L t s     0 �        p    ���    7���  &    v                      ���    /���  ;    l                    ���   ���� �   �         0            o��@  ?���� @  0     �   �             w��0  ���� 0  `    �  �         @   ����  ����@ �  �@     �  �      �  �   ����  r����   �  r�     x                ��������߀  x��         |             �����w����   �t       ��         p    ����������  ��      ���        ��    ��������}�@� ���  �     ?�         �     ���������     �                           =���������                                 ���������                               ���������                                  {�������x  �      �                       ���������         @                       ������{�  �     �                        ���������                                   ���������                                }�������                                   �������                                   �������   @                            �������                                                                   Q Q  g�����0   �8  �                         �?���}�   @�  �                      ~�����d   �    @�                        n������       D                        ��������                            ���������  H@    	                        ^�������`  �      B�  �     �             ���������  B      !          @            ���������            �      �            ���������       P                       ���������                            /���������                              [��������� $@                             �����������(        
 @�       �            �����������A        A                     m�������� �   �   $�                      _���0��� �   ��  �   �                ����  o���    p   @   ���               �����'�����H  �'�      �`              ��� @f�����  �O�      �              o���bF����  o�O��      �              ����J����  ��J��      `w�        #     ���p��_���  x���`     �p �       p     ���� ����  ����      p @             ����   W���@ ��X         �              �����L�����@ �泀�      ��P       �@�    �����G���� �3�D  @  ��8       ���    ��� �!���� ���b       `        @    �����7���� ���6     � �      � �   ���� ����  ,���     ��      � �    ���������  X��      ���      � �   ������
��  X�!�
�     ?=�~        |   ���?�~��  8?� ��    @>�>      >  >   �� >�>���  �? ~�    @|�ߟ      <     ���z@�/?��  �z�b�@    @}^�_�     x     ������?��  ���P�@    @z���      �    ��`����� p�    ����        �  ��@������ pX�    �������         �  ��@s���� `��    ��_�w��      �  �  ��@(�
��� `"�    �������         �  ��@X���� `"�    �������         �  ��@(�
��� `"�    �������         �  ��@S���� `��    ��_�w��      �  �  ��@�ǈ��� `	H�    �������         �  ��`����� `�    ����         �  �����Ѕ?��  ��P�@    @z���            ���zs����  �z���     @�\_��     x O   ��5��.����  �� .݀    [�����     �  �   ��������  /�  �    _�����     �  ?�   ���_�������  O_� ��     ?�}��       |�   ���������  O��c�     >����     � �~   ����������  %����     ���~      ��|   ����������� #�����     ��<      ��<   ���������� �����     ���8      ���8   �� �������� ����  @  ���8       ��   ����?� ����@ �>��      � 0       >�    ���@� ����@ `t�     �� `      p     ���   ���  0  `     �   �         @   ����  ����  �  �     �  �      �   �   ����  ����  �  ;�      x         `      o��Ӏ ������  S��       <               w���p�����  <|      � �             �����k����@  �l       ��         `    ����������   ��      ���        ��    ����O���߀   ���        ?�         �     �����������    �                           �����������                               ��������}�@�       �                       ���������                                  =���������                                 ���������                               ���������                                  {�������x  �      �                       ���������         @                       ������{�  �     �                        ���������                                   ���������                                }�������                                   �������                                   �������   @                            �������                                                                   Q Q    <�       � �       @                  �đ�      ;n        �                 >�>`      �� ��      @                  �����               @                ;��f     �l�      �                 L�?�_�     3��f      � @�               �������    @       �  �              g�����`    �   �     @                  ����?�   �   �`                        ;�����h   �    �                       �������                @              =�������                               [�������   $  ?�    @                  ��`?�v�  H��� �      �                n��  o��@  �   p D�  @  ���              }������`  � ��  �  ! �p B             ��'(p�� D ��/� @   �               ��� @�� @�H}�     �              ��0@_�� <
H`  � ��� �           
���@���  �@� P  � @            ���gv ��� 	 �ww �@   �              �� �z k�� 
@��z�l     s�        #"     +�� �� 7��  7 ���4    @ p       p     ;�   3�� �. ���2    p              W�    �� (�\ �                       W�P �L�
� ( � 泀
�@    ��       �@�   ��������	 ��3�  @ @ ���      ���   ��`� ����Bp����  �  `�       @ �  ��`����߀P`����   �� ��     � � �  ���� �_� R����` �� �� �     � � @  {�����_������@   ��� �     � � @  _�����_��!�@  ?=�~ �       | @  [��?�~ �����?� � �    >�> `     >  >    ���>�> �� �? ~ ��� |�ߟ p     <      �� z@�/ ��@�z�b� �  }^�_ p     x      �� ������H���P��    z�� 0      �    �� �� W��H  X    ����0          �� ��� _�� X@X	 H �����0           �� s� _��H�@X    �_�w�0      �    �� (�
 _��H"@X    �����0           ��X�@_�� "@X	 H �����0           ��(�
@_��H"@X    �����0           �� S� _��H�@X    �_�w�0      �    �� �ǈ _�� 	H@X	 H �����0           �� �� _��H  X    ����0           �� ��Ѐ���H	��P��    z�� 0            ��zs��@�z��  �\_ p     x O    ����.@�� ž .@������߀p    �      [�����������  ��   ������`    ��  ?�`  _��_������_� ��� ��}���    �  |��  {�}/���?����}��c���  �����    |� �?�  ��4w����� R 7����� ������?�    0���  ��������߀P������   ����     ���  ����������B������  �����     ����  ��� ������	 � ���� @ p ���       ��   W�L ?� >�� ( � >� ~ @  0 �        >�    W� � ?�� (�D t ~   8 �        p    ;�    /�� �"    n                    +��    o�� @    l                    ���   ��� 
 �   �         0            ��@  ���  `  �     �   `             ���  ���  �  �   @   @         @   ��  ��x  ��  =� �    �  �      �  �   ���  r���   ���     x                ��������   X�?�       ?  |             ����u���  ! 7�v B     ��         p    ��������  @ ��      ���        ��     ���������    ���        �         �      w�������   @ �                          /�������                                �������         @                         �������                                  �������                                   �������     @                             w�����@    �  �                          ~���      � @�                           /��o��      �                            �����       @                           �����      @                              ��o��       �                             ;���       @                                                          Q Q    <�       � �       @                  �đ�      ;n        �                 >�>`      �� ��      @                  �����               @                ;��f     �l�      �                 L�?�_�     3��f      � @�               �������    @       �  �              g�����`    �   �     @                  ����?�   �   �`                        ;�����h   �    �                       �������                @              =�������                               [�������   $        @                  ������v�  H�     �                        n������@  �  �  D�  @                   }��0��`  �  ��  �  !  �  B             ���  o�� D   p @    ���               �������� @ ��     �`              ��Ӏ ����  3�/�   � �  �            
��N@9��   �
Hy� P  0�             ���cF��� 	 �sG�@   @�             ��`�z_�� 
@p�z�`     �s� �       #"     +��������  �����    @ p `      p     ;��  ��� ������    p               W�    ��� (� � �                     W�� �L�g�� ( 7 泀d @   ��       �@�    ������3���	 .�3�2  @  ��       ���    ���� ����B L���   0  `        @   �������߀P X���     � �      � �    ��P� �
�� R ����
  ��  ��      � �   {��������� ����   @���      � �    _����� ��!�   @?=�~�       |   [�`?�~����`?� ��    �>�>�     >  > �  ��@>�>�� `? ~��� �|�ߟ�     <   �  ��@z@�/��@`z�b��  �}^�_�     x   �  ��@��󐂿��H`��P��    �z���      �  �  �����_��H�`    �����        @  �������� �X`	 H ������         @  ���s���H��`    �_�w��      �  @  ���(�
��H�"`    ������         @  ���X�_�� �"@	 H ������         @  ���(�
_��H�"@    ������         @  ���S���H��`    �_�w��      �  @  ����ǈ�� �	H`	 H ������         @  �������H �@    �����         @  ��@��Ђ���H`�P��    �z���          �  ��azs����@qz����  ��\_�     x O �  ��e��.ǿ�  e� .���� ����߁�    �  ��  [�o������� o�  ǀ    �������    �  ?À  _��_���� �_� ��   O�}���      }�   {�5������ ���c��   N����     � �   ��������� R _����  ��  ���      ��~   ���������߀P _�����     ��>      ��>   ����������B /�����   ���>      ���   ��� �������	 /����  @  ���<       ��   W�� ?� ��� (  >�� @   �        >�    W� � ��� (��t�    � 8      p    ;��   ��� �
�  �       p             +��`  O�� @`  P    �   �         @   ���  ��� 
 �  �     �  �      �   �   ��L  ?��  L  @      �  �      @      ��3� ���   �� �    |         0      ������x  � ,��  �      |             ����g���   �h      ��         `    ���p���   p        ���        p     ���������  !  O�  B      ?�         �     ���������  @  �                           ���������                                   w�������   @                             /�������                                �������         @                         �������                                  �������                                   �������     @                             w�����@    �  �                          ~���      � @�                           /��o��      �                            �����       @                           �����      @                              ��o��       �                             ;���       @                                                          Q Q    <�       � �       @                  �đ�      ;n        �                 >�>`      �� ��      @                  �����               @                ;��f     �l�      �                 L�?�_�     3��f      � @�               �������    @       �  �              g�����`    �   �     @                  ����?�   �   �`                        ;�����h   �    �                       �������                @              =�������                               [�������   $        @                  ������v�  H�     �                        n�������@  �      D�  @                   }�������`  �       �  !      B             �������� D      @                      ���0��� @  ��      �               ���  _���    `   �  ���  �            
����'����   �'�  P  �`              ����F���� 	  3�O� @   �             ����J��� 
@ o�J�      w�        #     +��X����   �����    @  p       p     ;�  ?�� �8���@    �p�             W�@  �� (�p�    �   �              W����L���� ( �況� @   ��`       �@�    ����������	 ��3��  @  ��p       ���    ���� �����B �����     `0        @   ������K�߀P ���L    � �8      � �   ���� �+�� R ���h  �� ��      � �   {�����5���� .��6    ���      � �   _������ ,�!�   ?=�~        |   [��?�~���� \?� �      >�>      >  >   ���>�>
��  X? ~ ��  |�ߟ      <     ���z@�/��@ Xz�b�    }^�_      x     ��Є�����H X��P�      z��       �    ��0����H ��    @����           �� �����  �X�	 H @�����            ���s����H ���    @�_�w�       �    ���(�
���H �"�    @�����            ���X����  �"�	 H @�����            ���(�
���H �"�    @�����            ���S����H ���    @�_�w�       �    ��0�ǈ��  �	H�	 H @�����            ��0����H ��    A����            ��[��Њ��H ۅP��    'z��G            ����s�����@ _�����   ?}\_b     x OB   �����.���  _� .� �� ?�����     �  �   [�������� _  �     ?�����     >  >�   _������� .߂ ��   ?}��       }�   {���������� /��c�~    ����     � �|   ��������� R ����  �� ���|     ��8   ��������߀P �����    ��8     ��8   ����������B �����   ���8     ���   �����������	 ����  @  ���p      ��    W���?���� ( �>�� @   � `      >� @   W�0�o�� (�0tp   �� �      p @   ;��  ��� ����    �  �      �  �   +���  2��� @�  r�     x                ��S� ��� 
  ���      <               ���p���   l|       � �             ����k���   �l     ��         `    ������x  � ��  �    ���        ��    ���������   ���       ?�         �     ���������    ?�                           ���������  !      B                        ���������  @                               ���������                                   w�������   @                             /�������                                �������         @                         �������                                  �������                                   �������     @                             w�����@    �  �                          ~���      � @�                           /��o��      �                            �����       @                           �����      @                              ��o��       �                             ;���       @                                                          Q Q    <�       � �       @                  �đ�      ;n        �                 >�>`      �� ��      @                  �����               @                ;��f     �l�      �                 L�?�_�     3��f      � @�               �������    @       �  �              g�����`    �   �     @                  ����?�   �   �`                        ;�����h   �    �                       �������                @              =�������                               [�������   $        @                  ������v�  H�     �                        n�������@  �      D�  @                   }�������`  �       �  !      B             �������� D      @                      ��������� @                            ��������   �    �       �            
��������    p   P   �               ���� ���� 	  � � @    ?�               ����"/��� 
@ �"�      �@              +�����K���   ���     @ p0       p     ;�� u��� � 7���     p              W��  ��� (� N�9     0                 W��0�L��� (  �泜� @   @��        �@�    ���a���?���	 q�3�@  @  ����       ���    ���A� ß���B a��à    �  `�        @�   �������_�߀P ����@    � ��      � �@   ����� ���� R Ͽ���  �� ��`      � �    {���������� ����    ���p      � �    _�����_� �!�X   ?=�~0        |   [��?�~W���� ?� �P     >�>8      >  >   ���>�>/��  ? ~( �� |�ߟ      <     ���z@�//��@ z�b�,   }^�_      x     ��������H ��P�     z��       �    ��������H      ����           ���������  ,X 	 H �����            ���s����H ,�     �_�w�       �    ���(�
���H ,"     �����            ���X����  ," 	 H �����            ���(�
���H ,"     �����            ���S����H ,�     �_�w�       �    ����ǈ���  ,	H 	 H �����            ��������H ,     ����            ����Л���H �P�     ���     �      ����s����@ ����   �\_�     � O   �����.���  � .� �� �����     �  �   [��������� �  �     �����     �  ?�   _������ ߂ ��   ?}��       }�   {��o�������� ��c��    ����     � ��   ���g����� R ����  �� ����     ���   ���G�����߀P g����    ����      ���   ���1�����B 1��Ơ    �����      ����   �����������	 ����  @  �����      ����   W��L?��� (  �>�� @   p�       @>�    W���&��� (� vt'     8�       0p    ;�ɀ ���� � )� �       <             +���p3��� @ p4      � �         0    ��������� 
  ���       ��       � �    ���p?���   p@        ���        p     ���������    O�       ?�         �     �������x  �  �   �                       ���������                                ���������                                 ���������  !      B                        ���������  @                               ���������                                   w�������   @                             /�������                                �������         @                         �������                                  �������                                   �������     @                             w�����@    �  �                          ~���      � @�                           /��o��      �                            �����       @                           �����      @                              ��o��       �                             ;���       @                                                          