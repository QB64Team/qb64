��j  聘�                 �    `                                          �    `                                          �    `                                          �    `                                          0   �    `                                     0   �    `                                     0   �    `                                     0   �    `                                         �    `                                         �    `                                         �    `                                         �    `                                     �����y�xsl�                                    �����y�xsl�                                    �����y�xsl�                                    �����y�xsl�                                    �m�6 `���cm�                                    �m�6 `���cm�                                    �m�6 `���cm�                                    �m�6 `���cm�                                                                                                                                           7����}��cm�                                                                                                                                                                                              6�`�Ͷ�cm�                                                                                                                                                                                             6m�6`�Ͷ�a͘                                                                                                                                                                                             ������}�x1��l                                                                                                                                                                                                        �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             �                                                                                                   �                                                                                                   7�                                                 `                                                 /�                                                                                                   /�                                                 0�                                                                                                   `@                                                 _�                                                 q�                                                 .                                                                                                     ��                                                 a�                                                 �@                                                 @�                                                 ��                                                 ��                                                 |`                                                ��                                                �                                               ���                                                �                                                 ��                                               ��                                               ��                                               ��                                                ��                                               ��x                                               ��                                               �a�                                               ��                                               ��                                               ��                                               �`                                               ��                                               ���                                              ���                                              �                                               ��                                              ����                                              ?��                                              ��                                               ���                                              ���x                                              ���                                              � a�                                              �g�                     0                        7���                                             o�g�                                              /�`                                             9��                     ,                        /���                    0                        0����                                                                   `                         ^��                    ^                        ����                    p                        1���                    .                        . �                                               ���                    ߀                       ���x                    a�                       ����                    �                        I  a�                    @�                        �@ g�                    ��                       �� �                    À                       �@ g�                    |                        d� `                   �                        o@ �                                           {� �                  �                        @ ��                   �                         �                     �                         � �                                           � ��                  �                         � �                  �                         @ �                                            � ��                  ��                        � �x                  �                        � ��                  �                         @  a�                  �                        �  g�                  ��                        �  �                  �                        �  g�                  �                            `                  �                        �  �                  �?�                       �  �                 ��                       �  ��                 ��                                             ��                       �  �                 ���                       x  ��                 ?��                       �  �                 �>                         �  �                  ��                       �  ��                 ���                      x  �x                 w���                      �  ��                 ��                        �   a�                 ?��                       �   g�                 7����                      �   �                 h?��                      �   g�                 /��                        H   `                 7���                       �   �                 /����                     �   �                0�����                     �   ��                 > �                       H                    ``~��                      z  ��                _����                      �������                q�~��                      ������                .�                       $   �                  (���                      {�����                �����                     ������x                a�����                     ������                �P  �                      $  �a�                @� ��                     ?��� '�                �� ���                     h   ���                �� ��                     ��� '�                |H  �                      �����`                ��  ���                     ?����	�                �  ��~                     o������               ��  ���                     ����	��               �H  �                        �                 z  �                     �����               ?�  ���                    7�������               �  ��                    ?�����               9$   �p                        ��                z   ���                        ��               ^   ���                    7������x               z   ���                    <    ��               $                        �����a�               =   �                    �������               o   �>                    �������               }   �                    �������                   ��                         `                =   ��                    @    �                o   �π                   �    �               }   ���                   @    ��                   p0                    �                    �   q��                   �                    7�   ��                   �    ��               >�   q��                   �    �               	                        @    �                �   ?�                   �    ��               7�   �|                   �    �x               >�   ?�                   �    ��               	    ��                   @     a�               @   ��                   �     g�               �   ��                   �     �               @   ��                   �     g�               �    0`                         `               @    1�                   �     1�               �    ?��                  �     o�              @    1��                  �     9��              �                             V               �    �                  �     2�              �    ��                  x     /��              �    �                  �     >�              @    �                    �     �               �    ��                  �     ��              �    �<                  x     7�x              �    ��                  �     ��              @     `�                   �     (a�              �     c�                   �     
g�              �     �                  �     �              �     c�                  �     g�                    0                   H     	`              �     �                   �     �              �     ��                 �     �             �     ��                 �     ��                                      H                   �     ?�                  z     �             x     ��                  �     ��             �     ?�                  �     �              �      �                   $     	�              �      ��                  z     
��             x      �<                  �     ��x             �      ��                  �     ��              �      0�                  $     �a�              �      3�                  =     g�             �      ?�                  o     ���             �      3�                  }     g�              H      0                       
��`              �      �                  =     �             �      ��                 o     ��            �      ��                 }     ���             H                             U              z      ?�                 �    �             �      ��                 7�    ���             �      ?�                 >�    ��             $       �                  	     U�              z       ��                 �     ���             �       �<                 7�    v�x             �       ��                 >�    ���             $       0�                 	      � a�             =       3�                 @    � g�             o       ?�                 �    v �             }       3�                 @    � g�                    0                 �     � `             =       �                 @    P �             o       ��                �    � �            }       ��                @    � ��                                    �     T              �      ?�                �    P �            7�      ��                �    � ��            >�      ?�                �    � �            	        �                 @     T �             �       ��                �     � ��            7�       �<                �     � �x            >�       ��                �     � ��            	        0�                @     (  a�            @       3�                �        g�            �       ?�                �     �  �            @       3�                �     p  g�            �       0                      �  `            @       �                �        �            �       ��               �        �           @       ��               �        ��           �                                            �       ?�               �        �           �       ��               x        ��           �       ?�               �        �           @        �                 �        �            �        ��               �        ��           �        �<               x        �x           �        ��               �        ��           @        0�                �         a�           �        3�                �         g�           �        ?�               �         �           �        3�               �         g�                    0                H         `           �        �                �         �           �        ��              �         �          �        ��              �         ��                                   H                    �        ?�               z         �          x        ��               �         ��          �        ?�               �         �           �         �                $         �           �         ��               z         ��          x         �<               �         �x          �         ��               �         ��           �         0�               $          a�           �         3�               =          g�          �         ?�               o          �          �         3�               }          g�           H         0                         `           �         �               =          �          �         ��              o          �         �         ��              }          ��          H                                             z         ?�              �         �          �         ��              7�         ��          �         ?�              >�         �          $          �               	          �           z          ��  @          �         ��          �          �<  @          7�         �x          �          ��  �          >�         ��          $          0�              	           a�          =          3����          @          g�          o          ?�  �          �          �          }          3����`          @          g�                    0���           �          `          =          �  �          @          �          o          ����P          �          �         }          ����          @          ��                                �                    �         >  `          �                    7�         ����           �          ��         >�         ?����          �          �         	           �             @          �          �          �  `          �          �          7�          ����           �          ��         >�          �����          �          ��         	                        @           a          @            `          �           f�         �          ���           �           �         @          ����          �           g�         �                                              @            �          �           �         �          ���P          �           ��        @          ���          �           ��        �                                               �           ���          �           ��        �          ���          x           ��        �          ���h          �           ��        @                          �                      �           � L          �           ��        �          � L          x           �x        �          � �          �           ��        @           H             �             �        �           � �           �           ��        �          � �          �           ��        �          �  �          �           ��                    H  �           H             `        �           � �           �           ��        �          � �          �           ��       �          � �          �           ���                   H �           H                     �           �            z           ��       x          � �           �           ���       �          �             �           ��        �           H              $             �        �           �  s           z           ���       x          �  �           �           ��x       �          �  N           �           ���        �           H  B           $             a�        �           �  �           =           �g�       �          �  n           o           ��       �          �  0           }           �g�        H           H                           `        �           �  s           =            �       �          �             o           ��      �          �  �           }           ���       H           H  `                                z           �  �           �           �       �          � �@          7�          ���       �          �   �          >�          ��       $           H              	             �        z           �  �          �           ��       �          �  <�          7�          ��x       �          �  �          >�          ���       $           H  �          	              a�       =           �  ;           @            g�       o          �  �          �          ?  �       }          �             @          ?  g�                  H             �             `       =           �  �          @            �       o          �  �          �          ?  �      }          �  8           @          ?  ��                 H             �                    �          �   �          �            �      7�         �  o�          �          ?  ��      >�         �              �          ?  �      	           H              @             �       �          �  0          �          >  ��      7�         �  0          �            �x      >�         �  �          �            ��      	           H             @              a�      @          �  �          �          <   g�      �         �  �          �          ~   �      @         �             �          ~   g�      �          H                            `      @          �  0          �          <   �      �         �  p          �          ~   �     @         �             �          ~   ��     �          H                                  �          �  0          �          <   �     �         �  �          x          ~   ��     �         �             �          ~   �     @          H               �              �      �          �  �          �              ��     �         �  �          x          ~   �x     �         �  8          �          ~   ��     @          H             �               a�     �          �  �           �              g�     �         �  �          �          �    �     �         �   �          �          �    g�                H   �           H               `     �          �  �           �               �     �         �  �          �         �    �    �         �  �          �             ��               H  �           H                    �          �              z               �    x         �  �           �         ƀ   ��    �         �              �         8�   �     �          H               $               �     �          �   4           z          8    ��    x         �  ~           �         ��   �x    �         �               �         D�   ��     �          H               $                a�     �          �   :           =          8     g�    �         �   �           o         ��    x     �         �   p           }         D�    g�     H          H   0                           �     �          �   Z           =          8     p    �         �   _           o         ��    �    �         �   0           }         D�    �     H          H                                     z          �              �                �     �         �   _           7�        ƀ    w     �         �   8           >�        8�    �     $          H              	                 p     z          �   -           �               �     �         �   /�          7�        �     �     �         �              >�             �     $          H              	                 �     =          �   �          @         @     �     o         �   ?�          �         �     �     }         �              @         �     �               H              �                �     =          �   �          @               �     o         �   �          �         �     ~�     }         �              @         �     �               H              �                �     �         �   �                    x     p�     7�        �   �          �         �    �w     >�        �   �          �         �    ��     	          H   �           @                p     �         �   �                     x    �p     7�        �   
8          �         �    ��     >�        �   �          �         �    ��     	          H                               p      @         �                       x    �      �        �             �         �    ��     @        �   �          �         �    ���     �         H                             �      @         �   ��                   x    ���     �        �             �         �   ���     @        �   ��        �         �   ���     �         H    �                            �         �   (                   x   ��      �        �   �        �         �   ?�      �        �   ��        �         �   ?��      @         H                             �p      �         �   � �                  x   ?�p      �        �           �         �  ���      �        �   ��        �         �  ��p      @         H                            �      �         �     y�                  <  ��      �        �   ?��        �         ~  ���      �        �   ���                 ~  ��                H     x�         �             8       �         �    ��                  <  �       �        �   �~�        �         ~  ~?�       �        �   ���        �         ~  �                 H    ��                    ��       �            ��         A         <  ��       x        �  ���        �         ~ ���       �        �  ���        W         ~ ���        �             ���        �                    �            � x�         ��        < ��        x        � ���        �        ~ ��        �        � �� �        ��        ~ ��         �            ���         	            p8         �         p � �          @@        8 �8        �        ������        ��        ���        �        ��� ��        V@        ���8         H           ���        ��          ��         �         �� ��          �    �  7����        �        ������        ��    G������        �        w�� ��        ��    �������         H          ���                �              z        �� �            �    ������          �        w���           �x   ����?��          �        �� �           �   ����?���          $          ���            ��          �p          {        � �             �   �  ~��p          �        w���            ���  �  ~?���          �        � �            ��   �  ~?��p          $          ��             H�        �          =�       ��              z���  �  ��          o�       w��             ��������������          }�       ��              z��?���?�����                   �              �2                     �        ��               �?���?����           7�       ��               ��?���?�����           >�       w�               ����������           	        h                 �@         �           �|   |  p                 ������������           ����������                 ��  �  ?��           ����������                 ������������                                     `���������            ���������                  c�?���?����                    �                 �?���?����            ����������                 c����������            ���������                                          |   |                    x?���?����            ����������                 �?���?����              |   |  �                 ���������            ���������                  �                                                �       �            ���������                  ����������              |   |                    �       �            ���������                   x?���?���              ��������                  ���������              ��������                   ���������             ��������                  �?���?����                                                                |   |                     �                      |   |                     �����                                            �                                                                        �                         ������                                                                   �                         ������                                                                    ��   �                    �                     ����                                            �    �                    �                                                                        �������                                                 �                                           ������@                                                                                              ~    �                                                 @                                            ~    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              � `�  ��                     |�                                                                                                                                                                           0    ��                     ��                                                                                                                                                                           0    ��                     ��                                                                                                                                                                           1�n�><�����                  ����ǜ�?�                                                                                                                                                                    1��lٻ��m�                  ��6l���ـ                                                                                                                                                                   1��lٳ>���m�                  �͛6o���߀                                                                                                                                                                   1��lٳf���m�                  �͛6l���                                                                                                                                                                    1��lٳf���m�                  �͛6l���ـ                                                                                                                                                                   1��f�3>���l�                  |���ǘ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                             