��]  |J� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         ����������������������������������������������������������������������������������������������������������������������������������������������������������������������� �                                       ������������������������������������������������������������������������������������������������������������������������������ ����������������������������������������������������������������������������������������������������������������������������������������������������������������������� �������������������������������������������                                       o���������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������             �                       p ���������������� ���������������������������������������������������������������������������������� ���������������������������             �    �                p ���������������� ��������������������������������������������������������������������������������� ��������������������������                  �8                p �����������������������������������������������������������������������������������������������������������������������������                  0 0                p �������������������������������������������������������������������������������������������������������������������������������                  p p                p �������������������������������������������������������������������������������������������������������������������������������                  `                  p �������������������������������������������������������������������������������������������������������������������������������                  �                  p �����������������������������������������������������������������������������������������������������������������������������                  �                  p ���������������������?����������������������������������������������������������������������������������?����������������������              �����              p ������������������� >g������������������������������������������������������������������������������ >g��������������������             ������              p ������������������� 3�`���������������������������������������������������������������������������� 3�`������������������             �0��3              p �����������������s����s����������������������������������������������������������������������������s����s��������������������             8>0�c              p ���������������������������������������������������������������������������������������������������������������������������             0<0 �              p �������������������������8����������������������������������������������������������������������������������8������������������             0x` 9�              p �����������������������1��������������������������������������������������������������������������������1������������������             `p� s�              p ����������������������C�������������������������������������������������������������������������������C������������������          ?� `�� �� ��           p �����������������?����� �����������������������������������������������������������������������?����� ���������������          ?� �8� �� ��           p ��������������������8� ��������������������������������������������������������������������������8� ���������������             �01�  �               p ���������������?��8�����x�������������������������������������������������������������������������?��8�����x�������������������            �0q�  �              p ���������������?ώ1�����q�������������������������������������������������������������������������?ώ1�����q�������������������            �0�  88              p ����������������c��������������������������������������������������������������������������������c�������������������������            �1��  0p              p ����������������<�������������������������������������������������������������������������������<������������������������            ��� 8 p�              p ����������������x�������������������������������������������������������������������������������x������������������������             �   �              p ���������������������������������������������������������������������������������������������������������������������������                                     p �������������������������������������������������������������������������������������������������������������������������������                                     p �������������������������������������������������������������������������������������������������������������������������������                                     p �������������������������������������������������������������������������������������������������������������������������������                                     p �������������������������������������������������������������������������������������������������������������������������������                                      p ���������������������������������������������������������������������������������������������������������������������������������������������������������������������p ��                                     ?�����������������������������������������������������������������������������������������������������������������������������p ��������������������������������������������������������������������������������������������������������������������������������������������������������������������p ������������������������������������������                                    ������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                �  �   �    � �p ������������������������������������������������������������������?������?�������������������������������������������������                
  ��         �p ���������������������������������������������������������������������������������������������������������������������������                
  ��         �p ���������������������������������������������������������������������������������������������������������������������������      ���        
q'��  � '0�p ������������������������������������������������lbq������������c1�����1������������������������������������������������������      �RQ        �	(��  Ȣ� ���p ������������������������������������������������o�������������}n���7]n����?_������������������������������������������������      S�_        y(��   ("� #��p �������������������������������������������������-�������������a`�����`�����_������������������������������������������������      4RP        �(��   ("�  ��p ������������������������������������������������˭�����������v�]o�����o�����_������������������������������������������������      4RQ        �Ȣ�  (�� @��p ������������������������������������������������˭�����������w7]n����]n�����_������������������������������������������������      �N        x��N  ��  @��p �������������������������������������������������-������������xa����8�q�����_������������������������������������������������                     �              �p ����������������������������������������������������������������������������������������������������������������������������                                   �p �����������������������������������������������������������������������������������������������������������������������������                                    �p ������������������������������������������������������������������������������������������������������������������������������������������������������������������p ��`                                    �����������������������������������������������������������������������������������������������������������������������������p ��������������������������������������������������������������������������������������������������������������������������������������������������������������������p ������������������������������������������                                    ������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p ��`                                    ����������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p ��`                                    ����������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p ��`                                    ����������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p ��`                                    ����������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p �����������������������������������������������������������������������������������������������������������������������������                                    �p ������������������������������������������������������������������������������������������������������������������������������������������������������������������p ��`                                    �����������������������������������������������������������������������������������������������������������������������������p ��������������������������������������������������������������������������������������������������������������������������������������������������������������������p �������������������������������������������                                    ����������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������         �      0                   p ������������������������������������������������������������������������������������������������������������������������������               0     �            p ������������������������������������������������������������������������������������������������������������������������������               0     �            p ������������������������������������������������������������������������������������������������������������������������������         �8�<��6<l�<���g�         p ������������������������������������������������������a��'�Ó���$��������������������������������������������������������         �3m���<fl�3f훶l�         p �����������������������������������������������������̒O�'Ù��g̙dI�?�������������������������������������������������������         ?0�>��8~l�0f͛6o�         p ��������������������������������������������������������?�3'ǁ��gϙ2dɐ?�������������������������������������������������������         0`f��<`l�0f͛6l          p �������������������������������������������������������矙3'ß��gϙ2dɓ��������������������������������������������������������         3m�f�p6f8�3f͛6��         p ������������������������������������������������������̒O�3�ə��g̙2d�?�������������������������������������������������������         8�>�`3<0�<��3�`        p ���������������������������������������������������������3�������3$�d�������������������������������������������������������                `  0                  p �������������������������������������������������������������������������������������������������������������������������������               �  �                  p �����������������������������������������������������������?������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p ���������������������������������������������������������������������������������������������������������������������������������������������������������������������� ��                                      ?����������������������������������������������������������������������������������������������������������������������������� ����������������������������������������������������������������������������������������������������������������������������������������������������������������������� �������������������������������������������                                       ��������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         ������������������������������������������������������������������������������������������������������������������������������