� �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 '''''''      '''''''''''''''    ''''''''''''            ''''''        '''''   '''     '''''''''''''     ''''   ''''''''''''''                                                                                                                                                '''''''     '''''''''''''''''    ''''''''''''''            '''''       '''''''  ''''    '''''''''''''''    ''''   ''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                '''''''''''''''''  ''              '''''''''''''     '''''''   '''         '''     ''''       '                                                                                                                                        '''''''''''''  ''''''''''''''''''   '''      ''      ''''''''''''''   '''   ''''''   '''      '''   ''''    ''''        ''                                                                                                                                       '''  '''''    '''       '''     '''''''   ''    ''''   '''       '''   '''    ''''       ''                                                                                                                                      '''  ''''    '''       ''    '''''''   '''      '''    '''       '''    '''    ''''       '''                                                                                                                                                     '''  '        ''   '''       '     '''     ''' ''      '''   '''      ''''   '''    '''       ''                                                                                                                                                     ''' ''        ''   ''' ''    ''''      ''' ''      '''   '''       '''   ''''    ''''      ''''                                                                                                                                                     '''''        ''   '''''''   ''''        '''' ''      '''   '''      ''''    '''    ''''    ''''                                                                                                                                                       ''''''''''        '''   ''''''''''''   ''''        ''' ''      '''    ''''''    '''    '''''''                                                                                                                                                       ''''''''''        ''   ''''''''''''''''    '''         '''''      '''    '''''''''''''    '''    '''''''                                                                                                                                                        ''''''''        ''    ''''''''''''''   ''''          ''''''''      '''    '''''''''''    ''''    '''''''''''''''                                                                                                                                                                 ''     '''''''''''''  ''''                 '''     '''''''''     '    ''''''''''''''                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     �����   ���� ����������� �������������             ����                                                                                                                                                                                                                                                                          ����   ���� ����������� ��������������           �����                                                                                                                                                                                                                                                                          ����  ����  ����        ����      ����          ������                  �������                                                                                                                                                                                                                     �������                                                                                           �����������                                                                                                                                                                                                                 �����������                    ��������                                         ����              ���������������                                                                                                                                                                                                             ���������������                  ��������   ��������    ��������������            ����             �����������������                                                                                                                                                                                                           �����������������                  ������    ��������    ��������������            ����            ������������������                                                                                                                                                                                                          ������������������                  ������    ����        ����   �����              ����            �������������������                                                                                                                                                                                                         �������������������                 ������    ����������� ����    �����             ����            �������������������                                                                                                                                                                                                         �������������������                  ����     ����������� ����     �����            ����            �������������������                                                                                                                                                                                                         �������������������                                                                                 �������������������                                                                                                                                                                                                         �������������������                                                                                 �������������������                                                                                                                                                                                                         �������������������                                                                                     �����������                                                                                                                                                                                                                 �����������                                                                                           �������                                                                                                                                                                                                                     �������                                                                                              �����                                                                                                                                                                                                                       �����                                                                                                ���                                                                                                                                                                                                                         ���                                                                                                 ���                                                                                                                                                                                                                         ���                                                                                                 ��                                                                                                                                                                                                                          ��                         ��������������   ������������    ������������    ����                     �      �                                                                                                                                                                                                                    �      �                 ���������������  ��������������  ��������������  �����                     �   ���                                                                                                                                                                                                                     �   ���                  ����       ����  ��������������  �������������� ������               �������������                                                                                                                                                                                                               �������������                                                                                        ������������                                                                                                                                                                                                                ������������                                   ����      ����  ����      ����   ����                � ��������                                                                                                                                                                                                                  � ��������                     ��������������  ����      ����  ����      ����   ����                 �      �                                                                                                                                                                                                                    �      �                     ��������������   ����      ����  ����      ����   ����                  �    �                                                                                                                                                                                                                      �    �                      ����             ����      ����  ����      ����   ����                   ����                                                                                                                                                                                                                        ����                       ���������������  ��������������  ��������������   ����                                                                                                                                                                                                                                                                          ���������������   ������������    ������������    ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �������������  �������������  �������������  �������������  �������������          �������������          �          ��  �������������  ��          �                                                                                                                                                                           ��          �  ��          �  ��             ��             ��                     ��          �          �          ��  ��             ��          �                                                                                                                                                                           �������������  �������������  �������������  �������������  �������������          �������������          ������������   �������������  �������������                                                                                                                                                                           �������������  �������������  �������������  �������������  �������������          �������������          ������������   �������������  �������������                                                                                                                                                                           ��             ��          �  ��                         �              �          ��          �          �          �   ��                   �                                                                                                                                                                                 ��             ��          �  �������������  �������������  �������������          ��          �          �          ��  �������������        �                                                                                                                                                                                 ��             ��          �  �������������  �������������  �������������          ��          �          �           �  �������������        �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         �                      �                                                                         �                                                 �                                                                                        �                                �                                    ����������  ���   �������� ���     ���   �������    ����������   ���������           ����������  ����������  ���   ��������         ����       ���             ���          ���������  ����������  ����������          ����������    ���������� ��      ���          ����������  ��      ���                                    ����������  ���  ��������  ���     ���  ���������   ����������   ����������          ���������   ����������  ���  ��������          ����      ����             ���          ���������  ����������  ���������           ����������   ����������  ���     ���          ����������  ���     ���                                    ���     ��� ��� ���        ���     ��� ���     ���  ���     ���  ���     ��          ���         ���     ��� ��� ���                �����    �����             ���         ���     ��� ���      �� ���                 ���     ��� ���          �����   ���          ���     ��� �����   ���                                    ���     ��� ��� ���        ����������� ���     ���  ���     ���  ���      ��         ���������   ���     ��� ��� ���                ������  ������             ���         ���     ��� ���     ��� ���������           �����������  ����������  ������  ���          ���     ��� ������  ���                                    ����������  ��� ���        ����������� �����������  ����������   ���      ��         ��������    ����������  ��� ���                ��� ��  �� ���             ���         ���     ��� ����������  ��������            ����������    ���������  ��� ��� ���          ����������  ��� ��� ���                                    ����������  ��� ���        ���     ��� �����������  ����������   ���      ��         ���         ����������  ��� ���                ��� �����  ���             ���         ���     ��� ���������   ���                 ���     ���           �� ���  ������          ����������  ���  ������                                    ���     ��� ��� ���        ���     ��� ���     ���  ���     ���  ���     ��          ���         ���     ��� ��� ���                ���  ����  ���             ���         ���     ��� ���         ���                 ���     ���          ��� ���   �����          ���     ��� ���   �����                                    ���     ��� ���  ��������� ���     ��� ���     ���  ���     ���  ����������          ����������  ���     ��� ���  ���������         ���   ��   ��� ���         ����������   ���������  ���         ����������          ����������    ���������  ���    ����          ���     ��� ���    ����                                    ���     ��� ���   �������  ���     ��� ���     ���  ���     ���  ���������           ���������   ���     ��� ���   �������          ���        ��� ���         ���������    ���������  ���         ���������           ����������   ����������  ���     ���          ���     ��� ���     ���                                              �                                      �            �                                            �                                     �                                       �                                                                                     �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ���������������         ��������   ����������   ����     ���  ���������������               ����   ����   ��������   ������  ������ �����������  �����������          ��������   ������������   ��������   �����   ���                                                                                                          ���������� ����        ����������  �����������   ���    ����  ���������� ����               ����   ����  ����������  ������  ������ ����������  �����������          ����������   ����������   ����������  ������  ���                                                                                                          ���������  ����       ������������ ������������  ����   ���   ���������  ����               ����   ���� ������������ �������������� ���������  �����������          ������������   ���������  ������������ ������� ���                                                                                                          ���������  ����       ����    ���� ����    ���    ���  ����   ����       ����               ����������� ����    ���� �������������� ����        ����������          ����    ����      ���     ����    ���� �����������                                                                                                          ���������  ����       ����    ���� ����������     ���� ���    ���������  ����               ����������� ����    ���� �������������� ���������   �����������         ����    ����      ���     ����    ���� �����������                                                                                                          ��������   ����       ����    ���� �����������     �������    ��������   ����               ����������� ����    ���� ���� ���� ���� ��������     ����������         ����    ����      ���     ����    ���� ���� ������                                                                                                          ����       ���������� ������������ ����    ����     �����     ���������� ����������         ����   ���� ������������ ���� ���� ���� ����������          ����        ������������      ���     ������������ ����  �����                                                                                                          ����       ����������  ����������  ����    ����     ����      ���������� ����������         ����   ����  ����������  ����  ��  ���� ����������  �����������          ����������       ���      ����������  ����    ���                                                                                                          ����       ���������    ��������   ����    ����      ���      ���������  ���������          ����   ����   ��������   ����      ���� ���������   ����������            ��������        ���       ��������   ����     ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �� ��       �����������  �� ��       �����������            ���������� ��      ��  �� ��        �� ���������� ����������  ��  ���    �� �������  ����������                                                                                                                                                                     �� ��       �����������  �� ��       �����������            ���������� ��      ��  �� ��        �� ���������� ����������  ��  ����   �� �������  ����������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     �� ��       ��       ��  �� ��       ��       ��            ���������� ����������  �� ��        �� ���������� ����������  ��  �� ��� �� ������   ����������                                                                                                                                                                     �� ��       ��       ��  �� ��       ��       ��            ���������� ����������  �� ��        �� ���������� ����������  ��  ��  ����� ������    ���������                                                                                                                                                                     �� �������� �����������  �� �������� �����������            ��         ��      ��  �� ��������  �� ��         ��          ��  ��  ����� �������� ����������                                                                                                                                                                     �� �������� �����������  �� �������� �����������  ��        ��         ��      ��  �� ��������  �� ��         ��          ��  ��   ���� �������� ����������                                                                                                                                                                                                                       ��                                                                                                                                                                                                                                                                                                                              ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   