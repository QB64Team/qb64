�`  �X�]                      �     6     0� �                                          �     6     0� �                                          �     6     0� �                                          �     6     0� �                                         3 � `     �0� �                                         3 � `     �0� �                                         3 � `     �0� �                                         3 � `     �0� �                                         0 � `     �0� �                                         0 � `     �0� �                                         0 � `     �0� �                                         0 � `     �0� �                                         0<�p<�6y�`9ͳ�<�8                                        0<�p<�6y�`9ͳ�<�8                                        0<�p<�6y�`9ͳ�<�8                                        0<�p<�6y�`9ͳ�<�8                                        fٳ`����m��c3fٰ                                        fٳ`����m��c3fٰ                                        fٳ`����m��c3fٰ                                        fٳ`����m��c3fٰ                                        ~߰`>��}��1���0fٰ                                        ~߰`>��}��1���0fٰ                                        ~߰`>��}��1���0fٰ                                        ~߰`>��}��1���0fٰ                                                                                                                                                                  `�0`f��͛���0fٰ                                                                                                                                                                                                                               3fٳ`f��͛`m�6l3fٰ                                                                                                                                                                                                                               <�0>�6}�08�3�<�3l                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ��      �`                                               ���      �p                                               ���      ���                                                 `       �                                                ?�      ���                                               ��      7���                                               ���      ���                                                ?�       ���                                               !��      /��                                               >?��      o��                                               ?���      ���                                               ��       ��                                                      ���                                               }��      _���                                               ?���      ?��                                               B        ��                                 �          =��     ���                         �        �          {���      ���            0            �        �          ?���     ?��                                   �          D         ?��           <            �       �          =��     ?���  0         <            �       �          w��      ?��  8         8            ��       �          ?����     ���           8             �        �          H         ?��           :            �        |�            �     ?���  6         9            ��       |�         ���      ?���  >         >            ��       ?��         ����     ���           8                    <�                  ?���  �        ;�           �        ���           �     ?���  3�        8�           7��       ���         w���      ?���  ?�        ?�           ?��       ��         ����     ���           8�                    s��                  ?���  �        ;�           ��      ���          ^ �     ?���  7�        8�           o��      ���         ���      ?���  ?�        ?�           ��       ���         ����     ���           8�            @       ���                   ?���  x        ;�           ?��      ��p          �{��     ?���  3�        8�           ���      ��p         ���      ?���  ?�        ?�           ���      ���         ����     ���           8�                    ��p                   ?���  �        ;�          ��      ���          �ߡ�     ?��_  7�        8�          ���      ���         ���      ?��c  ?�        ?�          ���      ���         ����     ���           8�           @        ���                   ?��   �       ;�@          ���      ��         o���     ?��  3��       8�@         ��      ��         ���      ?���  ?��       ?��         ���      ���         ����     ��           8�           �        ��                  ?��   ��       ;�         ��      ��         ���     ?��|  7��       8�         ���      ��         ���      ?���  ?��       ?��         ���      ���         ����     ��~           8�                    ��                   ?��   �       ;�         ���      ���          ��À     4|��  3��       8�         ���      ���         ���      4|�  ?��       ?��         ���      ���         ����     ��           8�                   ���                   4|    ��       ;�          ���      ���         ����     0&?�  7��       8�         ���      ���         ���      4��&  ?��       ?��         ���      ���         ����     {.?�           8�                    ���                   0     ��      ;� @        ���      ���         ���      0Y��  3���      8� @        ���      �F         ���      ?��  ?���      ?���        ���      ���         ���      p�           8�                   �@                   0     ���      ;�           ���      v,         ��^      RT��  7���      8�          ���      
���         ���      _���  ?���      ?���        ���      v<         ���      0  &           8�           [                                   ��      ;�           �_�      ��         ��<      _���  3���      8�          ���      �n�         ���      _���  ?���      ?���        �z�      �0         ���      0  L           8�                                                ���      ;�           ���      ���         ��x      _��X  7���      8�          ���      ���         ���      _��`  ?���      ?���        ���                 ���      0  �           8�                                                ��      ;�           ���      ���         ���      o���  3���      8�          ���      ���         ���      o���  ?���      ?���        ���      �         ���       0           8�                     �                          ���      ;�          ��      wj�         ���      o��`  7���      8�          ���      ��         ��       o���  ?���      ?���        ���       �j          ���       `           8�                     j                          ��      ;��@         ��      ��         ���      o���  3���      8ڠ@        ���      ��         ��       o��   ?���      ?���        ���       �           ���       �  �       8��                                                ��      ;��         ?��      ���         �ǀ      o���  7��      8��@        ���      ���         ��       o��   ?��      ?��        ���       @ @         ���       	�           8�                                                 ��      ;�           ��      ��p         ��       o��   3���      8�           ���      ��p         ��       o��   ?���      ?���         ���         �         ��                    8�                                                 ��       ;� �         ��      ���         ��       ��   7��       8� �         ��      ���         ��       ��   ?��       ?��          ��                 ��         &            8�                                                 �       ;�           ��       ���          �<       ��   3��       8� �         ?��       ���         ��       �0   ?��       ?��          ?��                 ��         �            8�                                                 ��       ;�           �        |�         A:x       �X   7��       8�           ��       |�         ��       �`   ?��       ?��          ��       �          ��        �            8�                                                                        ��       �          @��       �                          ��       �          ��       ��                          ��                   ��        0                                                                                               �           i�       ?�`                          �        �          �        ��                          �                    ?��        
`                                                @                                                             �       ?��                                                ?�        ?+                                                 ?��        ��                                                                                                             �       ��                                                �        f                                                 ��        ��                                                                                                                                                                     �                                                         �        �                                                                                                             �        �                                                                                                              �        �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          ��  �    0          �  �    ��          �      �                                                                                                                                                                                           �  ` �    1�          �  ��   ��          0      6                                                                                                                                                                                           �  ` �    00          �  ��   ��          0                                                                                                                                                                                                 �y�s��    0>s���      ��|珀   ��       3��>    �y�x                                                                                                                                                                                       ��fl�    0;fm�`      �v�ـ   ��3m�       �m�3f    lͶ�                                                                                                                                                                                       �}�g��    03fm��      ��f�ـ   ��3m�       �?f    lͶ�                                                                                                                                                                                       �ͳf�    03fm�       ��f��   ��3m�       m�0f    lͶ�                                                                                                                                                                                       �ͳfl�    1�fm�`      ��f�ـ   ��3m�       m�3f    6lͶ�                                                                                                                                                                                       �}�3��    3cͳ�      ��fg��    ��m�       홞>    �ly�x                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               �                                    @                                                                                                                                                                                                           �   c   �                �`� �   @           >                                                                                                                                                                                            �   c   �               � � �   @           3 �                                                                                                                                                                                            �   c   �               � � �   @           3 �                                                                                                                                                                                            �   c<�9���             ��o��<y�   @           3v���                                                                                                                                                                                           ����fͳm�6c����      �����nٳf�����      �����>fͷ`�����                                                                                                                                                                                           cf�?1�7�              ��lٳ`}�                3f��`                                                                                                                                                                                                cf�0�6               ��lٳ`̀                3f�f`                                                                                                                                                                                                cfͳm�6`              �slٳf̀                3fͶ`                                                                                                                                                                                                c<�9���               �clϳ<}�                >fl�`                                                                                                                                                                                                                        `                                                                                                                                                                                                                                                  �                                                                                             