�l  �z��                 `                                              `                                              `                                              `                                             �` 0                                           �` 0                                           �` 0                                           �` 0                                            ` 0                                            ` 0                                            ` 0                                            ` 0                                           g�8<��ny����<��<                               g�8<��ny����<��<                               g�8<��ny����<��<                               g�8<��ny����<��<                               3lٰf��l��m���f                               3lٰf��l��m���f                               3lٰf��l��m���f                               3lٰf��l��m���f                               �o�0f�������0>͛~                               �o�0f�������0>͛~                               �o�0f�������0>͛~                               �o�0f�������0>͛~                                                                                                                                       �l03f�����͛0f͛`                                                                                                                                                                                           �lٰ3f́�l͛m�0f͛f                                                                                                                                                                                           g�<���fy���0>��<�                                                                                                                                                                                                                                                                                                                                                                                                                           �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ?��                ��                ��                                                                                                                                                                       � |                �               | �                                                                                                                                                                      x  �             �                �  <                                                                                                                                                                     �   8                 �             8   �                                                                                                                                                                                     0                 �    `                                                                                                                                                                    0    �            �                                                                                                                                                                                         �     `                �                                                                                                                                                                                                          `           0     �                                                                                                                                                                                   0                 �      `                                                                                                                                                                                   @                                                                                                                                                                                                 �          �                                                                                                                                                                                         �       `                �                                                                                                                                                                                                          @                                                                                                                                                                                                                             �                                                                                                                                                                                                  @        @                                                                                                                                                                                                   �                                                                                                                                                                                          @                                                                                                                                                                                                   �        �                                                                                                                                                                                         @         @                                                                                                                                                                                                 �                           �                                                                                                                                                                                                         @                                                                                                                                                                                                                           �                                                                                                                                                                                                          �                                                                                                                                                                                              @          @                                                                                                                                                                                              �                                                                                                                                                                                      @                                                                                                                                                                                                      @                                                                                                                                                                                                 �      �                                                                                                                                                                                                �      �                                                                                                                                                                                    @           @                                                                                                                                                                                       @     @           @                                                                                                                                     @                                                   �     �                             �                                                                                                                    �            @                  @                        �                             �                                                                             @                  @                               @                  �                                                    @                                                                             @                  �                               �                  �                                                    @                                                                             �                  �                               �                                                                                         �                                                            �                                                                                                                                          �                                                                                                                                                                                                       �                                                                                                                                                  @                                       @            @                                                                                                @                                                 �                                       @            @                                                                                                �                                                                                        @            @                                                                                                                                                                                        @            @                                                                                                                                                                                          �                                                                                                                                                                                           �          �                                                                                                                          �                  �                             �                �          �                   @                 �                  �                               �                               `                 �                 �           `                �          �     �             �                 �                 �             `                  �                  �            P                 �                 �           X                �          �     �             �                 �                 �             @                 �                 �             �                 X                 �           �          @                    �           �                 �                 �             �                                   �            �                 �                 @           �          @     �               `           �                 ,                 �             �                                                �                 �                 .�           �          @     7<               .�           ��                �                 ,            �                                                O�                                 ]<           o�         @     ,               ]�           �0                ��                >s                                              0            �                n�                �           _�         @     o�              �           ��                �0                |��            �                                 8            
��                ^��               t?�          
��         @     ���             v��           3                ; �                �0            0                 �                p            <�                5��               ���          ��         @     ���             ���          p�               ~@3               � �                            0 0                � �           ??�              ���               ���          ���        @    ���             �?�          L0               r0�              ��3                            0                � 0           ��              z�?�              ���          -|��        @    s���            ���          � �               �0              �0�            �               `                �            *��               ����              O�?�         +?�        @    ����            o���         ��3              � �              �0            0               �  �                           ��              ��3�              .����         Z���        @    ��?�            .����         =  �             �  3              0  �                           �  0                 �          T<?�             ���              3�3�         �<��       @    ���            ��?�         9� 0             �  �             >L  3                          �                   0          1� ��             _`?�             =��         �� ��       @    ���           ?��         z   �             �  0             �  �         0   �                                           �� 3�             �` ��             ��?�        �� ?�       @    �� ��           ����        s   3             $   �             	P  0         !   0                �                         a� �             �� 3�             !� ��        i� �       @    7� ?�           ߀ ��        v�  �            �   3             (   �         `�                  0                 �         1� ?�            w� �             @ހ 3�        � ��           w� �       �     ߀ ?�         �  0             �   �             (   3          �                               @   0         "�  ��            � ?�            �/@ �        �  ��            K� ��      �     /� �         @   �                0                �         @   �                            �            @�  3�            �  ��            @ ?�        �  ?�            �  ��      �     � ��        @   3                 �                0        @@   0                �                        @z  �            �  3�            �  ��        ~  �            �  ?�      �     �  ��         �   �            �   3             
    �        @                 �   0                �        �z  ?�            �  �            �  3�        ~  ��           �  �      �     �  ?�         �   0            �   �            
    3        �                  �                   0        �=   ��             �  ?�           �  �        ?   ��           �  ��     @     �  � @       P    �            @   0                �       �    �             @                           =   3�           @ �   ��           �  ?�       ?   ?�           �   ��     @     �  ��@       P    3            @    �                0           0           @ @    �                       �  �           � z   3�            �   ��       �  �           ~   ?�     @     �   ��@       (    �            �    3            �    �                      �      0             �    �       �  ?�          � z   �          @ �   3�       �  ��           ~   �     @     �   ?�@       (    0            �    �           �    3                      �                @  �    0       @  ���           =  �?�         �  �  ��       �  ���           ?  ���            �  ���       ?��  �            P���             C���             �                         �  @           ���3�           =��� ��           ����?       ������           ?������            �������            0            P     �           @                0                �           @           �����           �����           ��� O       ������           ������            ������       
����              +����              ����         ����             ����             /���         ����            �����           ���        ������           ������           �����        
                  (                  �                                                           ���� @           ����            ?���        ������           ������           ?�����                                            P                                                          �                                 8       �     ������           ������           ?�����                                            P                                                          ������           �����             �����  �     ������           ������           �����        �                 
                  (             �                                               �                 �             @   �      @     �    @           �               �           �                 
                  (              �                               @                 �                 �             �   @      @      �    @           �               �           @                                                 @                               �              @  �              @  �                @             �    �      �     �               �           @                                              @  @              @                              @  z              �  �                �             ~    �      �     �               �            �                 �                 
           @                 �   �                           �  z              �  �                �            ~          @     �               �            �                 �                 
           �                 �   �                           �  =                 �                �            ?          @      �               �            P                 @                            �                   @                             =                 �                �            ?                 �          �     �             P                 @                                               @                             �                z                 �            �               ~          @     �   @         (                  �                 �                                                �            �                z            @    �            �               ~                 �   �         (                  �                 �                                          @     �            @                =            �     �            �               ?                  �   �                           P                 @                                         �     @            @                =                 �            �               ?   @             �                              P                 @                                              @            �                �                z       �     �                �  �             ~            
                  (                  �                                                           �                 �                 z       @     �  @             �               ~            
                  (                  �                                                             �                 @                 =             �  �        �     �               ?                                                P                                                            �            @    @                 =            �          @     �               ?                                                P                         @                                  �            �    �                 �           �                �          �     �            �                 
                  (             �            �                                   �            �    �                 �           �               �          @     � @          �                 
                  (              �            �                                    �                �                 @            �               �                 � �          @                                                 @                                           @    �                �                 @            �               � @              �           @                                            @    @                                           @    z                 �                 �       �     ~ `              ��              �            �                 �                 
         @                       �                          �    z                 �                 �             ~ �          �    �               �            �                 �                 
         �                       �                          �    =                  �                 �            ?           @     �               �            P                 @                          �                      @                              =                  �                 �            ?           0     �           �    �`            P                 @                                                @                               �                 z                 �            �                ~`           0    ��            (                  �                 �                                                  �             �                 z                 �        �    �                �               �             (                  �                 �                                                  �                               8                  �        0    �            �    >                 �                               P                 @                                                 @                                                  �                         0    8             �    �                               @                                                                                                                                  �   8                 �             8   �                                                                                                                                                                     x  �             �                �  <                                                                                                                                                                      � |                �               | �                                                                                                                                                                       ?��                ��                ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      � `�  ��         ̀`             �         0                                                                                                                                                              0    ��         l `�             0     0                                                                                                                                                                 0    ��          `�             0     0                                                                                                                                                                 1�n�><��;`<��<     �|�y�<��y�      ��͹��3π                                                                                                                                                            1��lٻ�����f     ͳv�Ͷf���      ͳ3m�m�7m�n�                                                                                                                                                            1��lٳ>����>͛~      m�f���~��͘      3?m��3�f6l�                                                                                                                                                            1��lٳf����f͛`      m�f���`�f͘      30m�3c6l�                                                                                                                                                            1��lٳf���`f͛f     m�f�ͶfͶ͘      �3m�m�6m�l�                                                                                                                                                            1��f�3>��30>��<     ͟f`y�<��y�      �m�͙�g3��                                                                                                                                                                                                                                                                                                                                                                                      �        >                                                                                 