�i  ,|��                       �       0  0                                             �       0  0                                             �       0  0                                             �       0  0                                            3 � `                                                    3 � `                                                    3 � `                                                    3 � `                                                    0 � `                                                    0 � `                                                    0 � `                                                    0 � `                                                    0<�p<x�<7�                                           0<�p<x�<7�                                           0<�p<x�<7�                                           0<�p<x�<7�                                           fٳ`�6f�ـ                                          fٳ`�6f�ـ                                          fٳ`�6f�ـ                                          fٳ`�6f�ـ                                          ~߰`>��6~1��                                          ~߰`>��6~1��                                          ~߰`>��6~1��                                          ~߰`>��6~1��                                                                                                                                                              `�0`f��6`3                                                                                                                                                                                                                         3fٳ`f͛6f��                                                                                                                                                                                                                        <�0>x��<7�6�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��            ��            ��            ��                                                                                                                                                                                       �"|           �"|           �"|           �"|          ݀            ݀            ݀            ݀          "             "             "             "                                                                    /���          /���          /���          /���        � \           � \           � \           � \                                                                                                                             c�"~0          c�"~0          c�"~0          c�"~0        ݁�          ݁�          ݁�          ݁�        "           "           "           "                                                                  �/���         �/���         �/���         �/���        A� \          A� \          A� \          A� \                                                                                                                           s���s�        s���s�        s���s�        s���s�      �  �         �  �         �  �         �  �                                                                                                           3��"�`        3��"�`        3��"�`        3��"�`      `݀1�        `݀1�        `݀1�        `݀1�       " @          " @          " @          " @                                                                 ����        ����        ����        ����       �� 8@         �� 8@         �� 8@         �� 8@       D          D          D          D                                                                �����|�       �����|�       �����|�       �����|�      f  �0        f  �0        f  �0        f  �0                                                                                                                         o�����v       o�����v       o�����v       o�����v      �0   `�        �0   `�        �0   `�        �0   `�        �D          �D          �D          �D                                                               ߿�����       ߿�����       ߿�����       ߿�����      @   &        @   &        @   &        @   &       �             �             �             �                                                                   ��������      ��������      ��������      ��������    C           C           C           C          �             �             �             �                                                                    >������{�      >������{�      >������{�      >������{�         �            �            �            �          �           �           �           �                                                              m��������      m��������      m��������      m��������         B@           B@           B@           B@                                                                                                                        ׿������X      ׿������X      ׿������X      ׿������X    (@     �      (@     �      (@     �      (@     �          !             !             !             !                                                              ��� ����     ��������     ��������     ��������    � �  @      �     @      �     @      �     @    @             @             @             @                                                                    ��� ���     ��������     ��������     ��������    �  x �        �             �             �           !             !             !             !                                                                    ���  ���     ���������     ���������     ���������   B �       B           B           B                                                                                                                             {��   ��     {��� ����     {��������     {��������    �   �      �  �        �            �                �            �            �            �                                                             ���   �~�    ���� ��~�    ��������~�    ��������~�   0   ` �       x �  �            �            �    �             �             �             �                                                                    ��    ��@    ���  ���@    ���������@    ���������@  	 �    D�    	 �   D�    	       D�    	       D�                                                                                                                      5��    ��`    5���   ��`    5���� ����`    5���������`  
      �    
    � �    
   �   �    
        �           @             @             @             @                                                            /��    ��    /���   ?��    /���� ���    /���������  @     @    @    @ @    @  8 �  @    @       @                                                                                                              [�     ��    [��   ���    [��  ����    [���������  $�    �	     $� `   0 	     $� �   	     $�       	                                                                                                                       ���     ?�X    ���    ��X    ����   ���X    ���������X  (      @ �    (  �     �    (       �    (   �    �  @�            @�            @�            @�                                                                    ���     ��    ���    ���    ����   ���    ����� ����  A        @    A      @    A     � @    A   <�  @                                                                                                             m��     ��   m��    ���   m���   ���   m���  ����  � @          �           �  0   `      �   �                @              @              @              @                                                           _��     ��   _��     ���   _���   ���   _���  ����  � @           �            �  @          �                                                                                                                     ��      ��   ���     ��   ���    ���   ����   ����  $ �          $      �     $  �         $                                                                                                                        ��      ��   ���     ?��   ���    ���   ����   ?���                 @                   �    @              @              @              @                                                                     ��      �~   ���     �~   ���    ��~   ����   ��~ @       �   @         �   @       �   @         �                                                                                                                 w�      ��   w��     ��   w��     ���   w���   ��� �           � @          �           �  @                                                                                                                           o�       ��   o��     ��   o��     ��   o��    ���  �           � @          �      �     �  �                                                                                                                      ��       ���  ��      ���  ���     ���  ���    ����           �               �             �              �              �              �                                                                     
��       ��  
��      ���  
���     ?���  
���    ����        �@           @          @ @           @                                                                                                                 
��       ��  
��      ���  
���     ���  
���    ����        �                                                                                                                                                            ��       ?��  ��      ���  ���     ���  ���     ����         @                                                                                                                                                       ��       ?��  ��      ���  ���     ���  ���     ����
        @   
           
  @         
          @              @              @              @                                                                     ��       ?��  ��      ���  ���     ���  ���     ���
@       @    
@           
@ @          
@      �                                                                                                                       ��       ��  ��       ���  ���     ���  ���     ���
@             
@           
@ @          
@      �                                                                                                                       ��       �@  ��       ��@  ��      ��@  ���     ?��@ @         �   @       �   @ �      �   @      @ �
              
              
              
                                                                      ��       ��  ��       ���  ��      ���  ���     ?���
             
           
  �         
       @   @              @              @              @                                                                     +�       ��  +�       ���  +�      ���  +��     ?����             �           � �          �      @                                                                                                                       +�       ��  +�       ��  +�      ���  +��     ?����@           �       �    �           �      @                                                                                                                       ?��       ��  ?��       ��  ?��      ���  ?���     ���  @       	@           �	@           	@             	@�             �             �             �                                                                     +�       ��  +�       ��  +�      ���  +��     ����@           �       �    �           �                                                                                                                               +�       ��  +�       ��  +�      ���  +��     ����@           �       �    �           �                                                                                                                               +�       ��  +�       ��  +�      ���  +��     ����@           �       �    �           �                                                                                                                               ?��       ��  ?��       ��  ?��      ���  ?���     ���  @       	@           �	@           	@             	@�             �             �             �                                                                     +�       ��  +�       ��  +�      ���  +��     ����@           �       �    �           �                                                                                                                               +�       ��  +�       ��  +�      ���  +��     ����@           �       �    �           �                                                                                                                               +�       ��  +�       ��  +�      ���  +��     ����@           �       �    �           �                                                                                                                               ?��       ��  ?��       ��  ?��      ���  ?���     ���  @       	@           �	@           	@             	@�             �             �             �                                                                     +�       ��  +�       ��  +�      ���  +��     ?����@           �       �    �           �      @                                                                                                                       +�       ��  +�       ���  +�      ���  +��     ?����             �           � �          �      @                                                                                                                       ��       ��  ��       ���  ��      ���  ���     ?���
             
           
  �         
       @   @              @              @              @                                                                     ��       �@  ��       ��@  ��      ��@  ���     ?��@ @         �   @       �   @ �      �   @      @ �
              
              
              
                                                                      ��       ��  ��       ���  ���     ���  ���     ���
@             
@           
@ @          
@      �                                                                                                                       ��       ?��  ��      ���  ���     ���  ���     ���
@       @    
@           
@ @          
@      �                                                                                                                       ��       ?��  ��      ���  ���     ���  ���     ����
        @   
           
  @         
          @              @              @              @                                                                     ��       ?��  ��      ���  ���     ���  ���     ����         @                                                                                                                                                       
��       ��  
��      ���  
���     ���  
���    ����        �                                                                                                                                                            
��       ��  
��      ���  
���     ?���  
���    ����        �@           @          @ @           @                                                                                                                 ��       ���  ��      ���  ���     ���  ���    ����           �               �             �              �              �              �                                                                     o�       ��   o��     ��   o��     ��   o��    ���  �           � @          �      �     �  �                                                                                                                      w�      ��   w��     ��   w��     ���   w���   ��� �           � @          �           �  @                                                                                                                           ��      �~   ���     �~   ���    ��~   ����   ��~ @       �   @         �   @       �   @         �                                                                                                                 ��      ��   ���     ?��   ���    ���   ����   ?���                 @                   �    @              @              @              @                                                                     ��      ��   ���     ��   ���    ���   ����   ����  $ �          $      �     $  �         $                                                                                                                        ]��     ��   ]��     ���   ]���   ���   ]���  ����  � @          �           �  @         �                                                                                                                            o��     ��   o��    ���   o���   ���   o���  ����  � @           �            �  0   `       �   �                                                                                                                           ���     ��    ���    ���    ����   ���    ����� ����  @         @    @       @    @     �  @    @   <�   @                                                                                                                      ��     ?��    ��    ���    ���   ����    ���������   �     @     � �         �          �  �                                                                                                                         ��     ��    ���   ���    ���  ����    ����������        �         `   0          �                                                                                                                                          ;��    ���    ;���   ?���    ;���� ����    ;����������                  @         8 �                                                                                                                                      /��    ��`    /���   ��`    /���� ����`    /���������`         �        �  �       �    �             �                                                                                                                      ��    ���    ���  ����    ����������    ����������     �             �                                                                                                                                                         ��   ���    ��� ����    ���������    ���������   � 0   `       �  x �        �             �                                                                                                                              ���   �}     ���� ���}     ��������}     ��������}      � �       �   �            �            �                                                                                                                       ���  ���     ���������     ���������     ���������      �                                                                                                                                                                        ���� ���     ���������     ���������     ���������    !  x �        !             !             !                                                                                                                              ���� ����     ���������     ���������     ���������    @  �         @             @             @                                                                                                                               ���������      ���������      ���������      ���������          !             !             !             !                                                                                                                         ��������      ��������      ��������      ��������                                                                                                                                                                                  7�������`      7�������`      7�������`      7�������`         �           �           �           �                                                                                                                        �������      �������      �������      �������     �             �             �             �                                                                                                                              ������       ������       ������       ������       �             �             �             �                                                                                                                             �����z       �����z       �����z       �����z        ��          ��          ��          ��                                                                                                                         �������       �������       �������       �������                                                                                                                                                                                    ^������        ^������        ^������        ^������      ! D@        ! D@        ! D@        ! D@                                                                                                                          ?������        ?������        ?������        ?������       " @          " @          " @          " @                                                                                                                           ������        ������        ������        ������                                                                                                                                                                    �����         �����         �����         �����                                                                                                                                                                                      }����          }����          }����          }����        "           "           "           "                                                                                                                             ����          ����          ����          ����                                                                                                                                                                                      ���           ���           ���           ���          "             "             "             "                                                                                                                               ��            ��            ��            ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           ?                        ?                                                                                                                                                                                                    0             3                          3                                                                                                                                                                                         0             0                          3                                                                                                                                                                                         >���          0���          ���          3���                                                                                                                                                                                      3훰          >훰          훰          훰                                                                                                                                                                                      ̓0          3̓0          ̓0          3̓0                                                                                                                                                                                      ̓0          3̓0          ̓0          3̓0                                                                                                                                                                                      3͛0          3͛0          ͛0          3͛0                                                                                                                                                                                      ��0          ��0          ��0          ��0                                                              