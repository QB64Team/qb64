��]  |J� ������������������������������������������������������������������������������������������������������������������������������                                          �                                        @�                                        @�                                        @                                          �                                        @�                                        @�                                        @                                          �                                        @�                                        @�                                        @                                          �                                        @�                                        @�                                        @                                          �                                        @�                                        @�                                        @                                          �����������������������������������������@�                                        @�����������������������������������������@���������������������������������������� �                                       @�                                        @�                                       @                                        �����������������������������������������@�                                        @�����������������������������������������@���������������������������������������� ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                      P@�                                        @��                                      P@�                                      P ��                                �    P@�                                 �     @��                                �    P@�                                      P ��                                �    P@�                                 �     @��                                �    P@�                                      P ��                              � �    P@�                               � �     @��                              � �    P@�                                      P ��                            � ?�    P@�                             � ?�     @��                            � ?�    P@�                                      P ��           >    >            � �    P@�            >    >            � �     @��           >    >            � �    P@�                                      P ��           >    >            � |    P@�            >    >            � |     @��           >    >            � |    P@�                                      P ��           |    |            � �<    P@�            |    |            � �<     @��           |    |            � �<    P@�                                      P ��           |    |            � �<    P@�            |    |            � �<     @��           |    |            � �<    P@�                                      P ��           �    �            ��<    P@�            �    �            ��<     @��           �    �            ��<    P@�                                      P ��           x    x            ��<    P@�            x    x            ��<     @��           x    x            ��<    P@�                                      P ��                           ��    P@�                            ��     @��                           ��    P@�                                      P ��                             ��    P@�                              ��     @��                             ��    P@�                                      P ��                  �          �     P@�                              �      @��                  �          �     P@�                  �                  P ��                  0          �     P@�                   �          �      @��                  �          �     P@�                  �                  P ��                 �0@         �     P@�                  ��         �      @��                 ���         �     P@�                 ���                 P ��       �        	�        > �     P@�        �        ���        > �      @��       �        ���        > �     P@�                 ���                 P ��      �     �  +\�        <��     P@�       �     �  ���        <��      @��      �     �  ���        <��     P@�                 ���                 P ��     @�  �� m�    � |��     P@�      @�  �� ���    � |��      @��     @�  �� ?���    � |��     P@�                 ?���                 P ��     ��� �?� a��J   �� x��     P@�      ��� �?� ���   �� x��      @��     ��� �?� ���   �� x��     P@�                 ���                 P ��     �?����  ��e   �� x��     P@�      �?���� ���   �� x��      @��     �?���� �����  �� x��     P@�                 �����                P ��    ������ �w�@�  �� ��      P@�     ������ _���   �� ��       @��    �����������  �� ��      P@�                �����                P ��    ����������h�  ?�� � |      P@�     �������� ����   ?�� � |       @��    �������������  ?�� � |      P@�                �����                P ��    �����>���>D����  ���� �      P@�     �����>���> ����   ���� �       @��    �����>���>�����  ���� �      P@�                �����                P ��    ���� <��<���� ���� �      P@�     ���� <��<����  ���� �       @��    ���� <��<����� ���� �      P@�                �����                P ��    ��� |�� |����p ���� �      P@�     ��� |�� |���� ���� �       @��    ��� |�� |����� ���� �      P@�                �����                P ��                ��p                P@�                 �����                 @��    ߟ� x� x����� �����      P@�                �����                P ��                ���x                P@�                 �����                 @��    �?> �� ������ �����      P@�                �����                P ��                ���8                P@�                 �����                 @��    �~| ��> ������ ����      P@�                �����                P ��                9��8                P@�                 �����                 @��    �>�|��<������ ?� ��      P@�                �����                P ��                y���                P@�                  ����@                 @��    �?����|������ ~� ��      P@�                �����                P ��                ����                P@�                 ���@                 @��    ?�����|������ �� ��      P@�                �����                P ��                %/���                P@�                  ���@                 @��    ?����?����������  �      P@�                �����                P ��                1fR$                P@�                   ���                 @��    �����?���������� < �      P@�                �����                P ��    �������A!���� <        P@�                   ?��                  @��    �������������� <        P@�                �����                P ��    ������$ ����x |        P@�                  #���                  @��    ������������x |        P@�                �����                P ��    �������  ��?x x> >       P@�                  ���                  @��    �������������?x x> >       P@�                �����                P ��   ��� �� �@ì�>x �< >       P@�                  r��<@                 @��   ��� �� ������>x �< >       P@�                �����                P ��   ����� �@��~� �< |       P@�                  u��                  @��   ����� ������~� �< |       P@�                �����                P ��   ����� � ��~��| |       P@�                  r��                  @��   ����� ������~��| |       P@�                �����                P ��   ����� ��;�� ���x �       P@�                  _�                  @��   ����� ����� ���x �       P@�                �����                P ��   �� >��> �s������x �       P@�                   @                   @��   �� >��> ��������x �       P@�                �����                P ��   �� <��< ����������       P@�                    "                   @��   �� <��< ����������       P@�                �����                P ��   �� |� | ����������       P@�    �� |� |   @  �����        @��                �����                P@�                �����                P ��   � > x� x �������? ��       P@�    � > x� x      ��? ��        @��                �����                P@�                �����                P ��     < �� �  �����x���       P@�      < �� �       �x���        @��                �����                P@�                �����                P ��     | ��> �  O���������       P@�      | ��> �       �����        @��                �����                P@�                �����                P �     |  >  c���@��?�  �       P �     |  >        ��?�  �       P �                 �����                 @�                �����                P �       x    <    �w���?�  �       P �       x    <         ��?�  �       P �                  �����                 @�                 �����                P �               A�~z ���  �       P �                    ���  �       P �                  ���                  @�                 ���                 P �                  �h  �            P �                       �            P �                  ?���                  @�                 ?���                 P �                    �            P �                       �            P �                  ���                  @�                 ���                 P �                    �  �            P �                       �            P �                  ���                  @�                 ���                 P �                    ��    >        P �                     ��    >        P �                  ���                  @�                 ���                 P �                     �             P �                     �             P �                   �                   @�                  �                  P �                     �             P �                     �             P �                   �                   @�                  �                  P �                     �              P �                     �              P �                                        @�                                      P �                     �>              P �                     �>              P �                                        @�                                      P �                     �|              P �                     �|              P �                                        @�                                      P �                     ��              P �                     ��              P �                                        @�                                      P �                     ��              P �                     ��              P �                                        @�                                      P �                     ��              P �                     ��              P �                                        @�                                      P �                      ��              P �                      ��              P �                                        @�                                      P �                      �              P �                      �              P �                                        @�                                      P �                                     P �                                     P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P �                                      P �                                      P �                                        @�                                      P ���������������������������������������� ���������������������������������������� �                                        @����������������������������������������                                                                                 �                                        @                                        ���������������������������������������� ���������������������������������������� �                                        @����������������������������������������                                                                                     �                                        @                                                                                                                              �                                        @                                                                                                                              �                                        @                                                                                                                              �                                        @                                                                                                                              �                                        @                                                                                                                              ������������������������������������������                                          