��]  |J� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         ����������������������������������������������������������������������������������������������������������������������������������������������������������������������� �                                       ������������������������������������������������������������������������������������������������������������������������������ ����������������������������������������������������������������������������������������������������������������������������������������������������������������������� �������������������������������������������                                       o���������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                               ����� p �������������������������������������������������������������������������������������������������������������������������������                               ����� p ����������������������������������    ����������������������������������������������������������������������������������������                               ����� p ����������������������������������    ����������������������������������������������������������������������������������������                               ����� p ����������������������������������    ����������������������������������������������������������������������������������������                            ����� p ����������������������������������    ����������������������������������������������������������������������������������������           p                ����� p ����������������������������������    ����������������������������������������������������������������������������������������           `                ����� p ����������������������������������    ����������������������������������������������������������������������������������������     8     8 �                ����� p ���������������������������������    ������������������������������������������������������������������������������������� 8    0�    0�                 ����� p ��������������������������������    ���������������������������������������?���������������������������������������?������ 0    �    �                 ����� p ��������������������������������    �������������������������������������  �������������������������������������  ������ 0   ��   ��                 ����� p �������� ?���� ?������������������    �������������������������������������  ������������ ?���� ?�������������������  ������ `����!���� ?            ����� p ����>�|����|��~|���������������    �������������������������������������  ��������>�|����|��~|����������������  ������ `����������ρ��           ����� p ����? ??�q�??�p>0~ ������������    �������������������������������������  ��������? ??�q�??�p>0~ �������������  ������ �σ������c���           ����� p ���0|>?���>?��`�>������������    �������������������������������������  �������0|>?���>?��`�>�������������  ������ ��������8cw            ����� p ���>Dp�~�x��>�ǜ����������������    ���������������������������������������?�������>Dp�~�x��>�ǜ�������������������?������ ����1��pg�8?            ����� p ���<��|����|����������������    ����������������������������������������������<��|����|��������������������������� 8`� `g�8            ����� p ���<������ǟ|��1���������������    �����������������������������������������������<������ǟ|��1����������������������������<x��ǌ             ����� p ���|9��������?8s���������������    �����������������������������������������������|9��������?8s����������������������������8�����            ����� p ���xq�����?���?0���������������    �����������������������������������������������xq�����?���?0������������������������� |<p�<�� �            ����� p ��������Ï����?1���������������    ����������������������������������������������������Ï����?1���������������������������p��9��8            ����� p ������q�����~a����������������    ��������������������������������������������������q�����~a����������������������������`;� �1��0�            ����� p �����y�?����?�|c� �������������������������������������������������������    ��������y�?����?�|c� ������������������������8���7��q�8q�                   p �����������xǎ��������������������������������������������������������������������������xǎ������������������������1� �<� a�0c�8                   p �����?���?�<����qϜ��������������������������������������������������������������������?���?�<����qϜ������������������������8q���x�� ��p��                   p ���ǎ��?�>���������������������������������������������������������������������ǎ��?�>��������������������������� �� �!�� @� A��                   p ����� ���~���߾ ?������������������������������������������������������������������� ���~���߾ ?�����������������������   �            �                    p ������������������ ��������������������������������������������������������������������������������� ������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p ��������������������������������������������������������������������������������������������������������������������������������  �         @   �           p ���_��}������������������������������������_��}�������������������������������������_��}������������������������������������   �  @�         �             p ����������o��������������������������������������o���������������������������������������o�������������������������������   �  @�         �             p ����������o��������������������������������������o���������������������������������������o�������������������������������,p�q�`�89��L�2�@r����'��9$   p ���ӏ��3�)���'���M��}58�8�������������ӏ��3�)���'���M��}58�8��������������ӏ��3�)���'���M��}58�8�������������2�"��(@�D%R	Jʀ
�+(�(��@�E$   p ����w�uu��f�������5�|��|�W[��}����������w�uu��f�������5�|��|�W[��}�����������w�uu��f�������5�|��|�W[��}���������"�"��@�|=%�H	"� z�*/�(��@�}T   p �����u��n��������t��}��}�Po�������������u��n��������t��}��}�Po��������������u��n��������t��}��}�Po�����������"�"��@�@E% D	����*((�AAT   p �����u}��n��������uu}����W���������������u}��n��������uu}����W����������������u}��n��������uu}����W�������������"�"��(@�DE%R	J�@��*(�(��A�D�   p ����w�uu��n������u�u}��}�W[��}�w��������w�uu��n������u�u}��}�W[��}�w���������w�uu��n������u�u}��}�W[��}�w�������"p�q�@Q8=$�L�2� z�*'''@�8�   p ���ݏ��;��������u߅}���������w�������ݏ��;��������u߅}���������w��������ݏ��;��������u߅}���������w�������                                    p �������������������������������������������������������������������������������������������������������������������������������                                    p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������        A                 �   p ������������������������������������}����������������������������������������}�����������������������������������������}������� @       A       �      �      p �����������������������������o���������������������������������������o����������������������������������������o������������� @       A       �      �      p �����������������������������o���������������������������������������o����������������������������������������o�������������l�0`x�y8&8��,��<r� r��8z��p  p ����q�㟇������8�8�&7Í8ߍ?)��3�a��������q�㟇������8�8�&7Í8ߍ?)��3�a���������q�㟇������8�8�&7Í8ߍ?)��3�a�������	IH�E�ED)D(�(��("(�� �D�(��  p �������o��Z���ֻ��}�Mm����_t�f��t��]w����������o��Z���ֻ��}�Mm����_t�f��t��]w�����������o��Z���ֻ��}�Mm����_t�f��t��]w������I @EE|$|/���("z/�� �|�(��  p �������Ὼ��ۃ��}�]m�݅�_u�n��u��]����������Ὼ��ۃ��}�]m�݅�_u�n��u��]�����������Ὼ��ۃ��}�]m�݅�_u�n��u��]������I" E	E@"@(��("�( � �@�(��  p ��������ߺ�����ݿ����]m��u��u�n��u��]�����������ߺ�����ݿ����]m��u��u�n��u��]������������ߺ�����ݿ����]m��u��u�n��u��]������	I�H"�E�ED)D(�(��("�(�� �D�(��  p �����n��o��Z���ֻ��}�]m��u�_u�n��u��]w��������n��o��Z���ֻ��}�]m��u�_u�n��u��]w���������n��o��Z���ֻ��}�]m��u�_u�n��u��]w������(�N0`x�y9�8
'�"Q�<z' r Q8z$�p  p ������ះ���9����8ݮ7Å�ߍ߮����a����������ះ���9����8ݮ7Å�ߍ߮����a�����������ះ���9����8ݮ7Å�ߍ߮����a�������       @                             p �������������������������������������������������������������������������������������������������������������������������������       @                       �      p ����������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                �  >�         p �������������������������������������������������������������������������������������������������������������������������  H      �        �       H     p ���߷�������������������������߷����������߷�������������������������߷�����������߷�������������������������߷����������  H      �        �       H     p ���߷�������������������������߷����������߷�������������������������߷�����������߷�������������������������߷����������0k9�r������c�8��� �08�0k,zp p ���ϔ���c�?1�k
p��m��N3?�L��
�ϔ��Ӆ������ϔ���c�?1�k
p��m��N3?�L��
�ϔ��Ӆ�������ϔ���c�?1�k
p��m��N3?�L��
�ϔ��Ӆ�������L�	E"� � U@Q�TD�) <���L� ��� p ���_�]���t�n�����o���5���[_���_�]�Muw�����_�]���t�n�����o���5���[_���_�]�Muw������_�]���t�n�����o���5���[_���_�]�Muw������H�A>� ��@�Q��|�(� � = H���� p ���_�A����n�*���l'��u��]����߷A�]u�����_�A����n�*���l'��u��]����߷A�]u������_�A����n�*���l'��u��]����߷A�]u������H�A � �UAQ�T@�(@ � E H���� p ���_�_���}�n�����k���u׿�^ߺ��߷_�]u�����_�_���}�n�����k���u׿�^ߺ��߷_�]u������_�_���}�n�����k���u׿�^ߺ��߷_�]u������H�	E"� �UAQ�RD�)  ��E4�H���� p ���_�]���u�n�����k���u���[_���_�]�]uw�����_�]���u�n�����k���u���[_���_�]�]uw������_�]���u�n�����k���u���[_���_�]�]uw����� (�9r N��@�O��8��� �<��(��zp p �����c���߱�+���l.��v;7�\��,��c�]���������c���߱�+���l.��v;7�\��,��c�]����������c���߱�+���l.��v;7�\��,��c�]�������                                   p �������������������������������������������������������������������������������������������������������������������������������           �                     �  p �������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������          �A��     
     ��  p ������������������a��}�������������_���������������������a��}�������������_����������������������a��}�������������_������  H   �     � �A        �  ��  p ���߷���o�����o���^��������������o��������߷���o�����o���^��������������o���������߷���o�����o���^��������������o��������  H   �     � �A        �  ��  p ���߷���o�����o���_��������������o��������߷���o�����o���_��������������o���������߷���o�����o���_��������������o��������0k"��2���8�A 2�s (���r@r��8��� p ���ϔ���&3��N)���_���a���f~5���?)��Xc?�����ϔ���&3��N)���_���a���f~5���?)��Xc?������ϔ���&3��N)���_���a���f~5���?)��Xc?������L���(J� �D��A�J�� (�*��� �D��� p ���_�]�]m��5�f��kX��]u��Z��ut�f��W]�����_�]�]m��5�f��kX��]u��Z��ut�f��W]������_�]�]m��5�f��kX��]u��Z��ut�f��W]������H����"� �|��A "�� (�
� � �|��� p ���_�A�]l��u�n��m^���]��n��|�u�n��WA�����_�A�]l��u�n��m^���]��n��|�u�n��WA������_�A�]l��u�n��m^���]��n��|�u�n��WA������H���� �@��A ��(�
��� �@��� p ���_�_�]m���u�n��n^���]}��v��}u�n��W_�����_�_�]m���u�n��n^���]}��v��}u�n��W_������_�_�]m���u�n��n^���]}��v��}u�n��W_������H���(J� �DQ�A J��)�*�@� �D��� p ���_�]�Ym��u�n��\���]u��Z��u�u�n��W]�����_�]�Ym��u�n��\���]u��Z��u�u�n��W]������_�]�Ym��u�n��\���]u��Z��u�u�n��W]����� (�I�2��Q8P�}�2�r@Ƙ��r r Q8��� p �����c��7��v���b��a��9g~5�ߍ߮��Xc�������c��7��v���b��a��9g~5�ߍ߮��Xc��������c��7��v���b��a��9g~5�ߍ߮��Xc�����                                     p �������������������������������������������������������������������������������������������������������������������������������         �                          p �������������?����������������������������������������?�����������������������������������������?������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������           8               �  p �������������������������������������_����������������������������������������_�����������������������������������������_������           D	             �  p ����������������������������������������������������������������������������������������������������������������������������           @	             �  p ����������������������������������������������������������������������������������������������������������������������������,x�<�0<䕀@�c��q�sNE��9�āǨ� p ���Ӈ�1���C���j��0�����~i�|;~8Wg�����Ӈ�1���C���j��0�����~i�|;~8Wg������Ӈ�1���C���j��0�����~i�|;~8Wg����� ��"�D��E�@9	�A(�� �QEYE$�(�� p ���Mw�~���]�_��i����k��]u�u���������W[�����Mw�~���]�_��i����k��]u�u���������W[������Mw�~���]�_��i����k��]u�u���������W[�������"�D��ET@�	���� �QEE$�訑�p ���]w�p���]�_�꫿���?wA�u�������~Wn����]w�p���]�_�꫿���?wA�u�������~Wn�����]w�p���]�_�꫿���?wA�u�������~Wn������"�D��ET@	 H�� �QE �E$�(�� p ���]w�n���]�_�꫿������_}�u����n���}�Ww�����]w�n���]�_�꫿������_}�u����n���}�Ww������]w�n���]�_�꫿������_}�u����n���}�Ww�������"�D	��E$@E	A(�� ��MQE#(�� p ���]w�n���]�_��ۿ�����]u�u�n��������V[�����]w�n���]�_��ۿ�����]u�u�n��������V[������]w�n���]�_��ۿ�����]u�u�n��������V[������x�<� <�$P8���q�r5�8��禘 p ���]��p���C���ۯ���0������n�|=�Yg�����]��p���C���ۯ���0������n�|=�Yg������]��p���C���ۯ���0������n�|=�Yg�����                                  p �������������������������������������������������������������������������������������������������������������������������������     x                             p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������   �|y��          (���       p ��������a���}����������������oA����������������a���}����������������oA�����������������a���}����������������oA�����������  H !B�    H        �P�        p ��������޽z����������������_���w�����������������޽z����������������_���w������������������޽z����������������_���w������������  H !B�    H         P�        p ��������޽~��������������������w�����������������޽~��������������������w������������������޽~��������������������w������������X�k!B� 2�s`k9��I8�)�P�        p ������޽~��a�������'��o��6��w���������������޽~��a�������'��o��6��w����������������޽~��a�������'��o��6��w������������	eL�!|��J���L�	%I�**��        p �����]�ރ~�]u�o�]�����o����ow��������������]�ރ~�]u�o�]�����o����ow���������������]�ރ~�]u�o�]�����o����ow������������	EH�!B� "��H�=%�U<�*�        p �����A�޽~��]��A�����o�����w��������������A�޽~��]��A�����o�����w���������������A�޽~��]��A�����o�����w������������	EH�!B� ��H�E% UD�*
�        p �����_�޽~��]}��_������o�����w��������������_�޽~��]}��_������o�����w���������������_�޽~��]}��_������o�����w������������	EH�!B� J��H�	E%"D`�)�        p �����]�޽z��]u��]����ݻ��U���w��������������]�޽z��]u��]����ݻ��U���w���������������]�޽z��]u��]����ݻ��U���w������������D�(�By�2�r(�=$�"<D)Ȉ"       p �����c�὆�a����c����û��7w����������������c�὆�a����c����û��7w�����������������c�὆�a����c����û��7w��������������                      @              p ������������������������������������������������������������������������������������������������������������������������������� �                   �              p �������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������O>�@  @  ( * @  @      � H      p �����������������������������_���������������������������������������_����������������������������������������_�������������P��
@  @  ( 
 @  @      �      p ���w������������������������_�������������w������������������������_��������������w������������������������_�������������P���@  @  ( 
 @  @      �      p ���w�u����������������������_�������������w�u����������������������_��������������w�u����������������������_�������������
P���X�OX��($�NI�IX9���X,�g�8� p ����w}�t����8�8��U����1����D�[��?�q�������w}�t����8�8��U����1����D�[��?�q��������w}�t����8�8��U����1����D�[��?�q������
P��JeQd(� �$�	QIQIdE$���P) �QE p ����w���뮛��}�W�U���������}[���k���������w���뮛��}�W�U���������}[���k����������w���뮛��}�W�U���������}[���k��������	P��JEQD/�'�*�QUQUDE$���P(�D_} p ����w���뮻��}�W�U���������a[������������w���뮻��}�W�U���������a[�������������w���뮻��}�W�U���������a[�����������Ј��EQD((�*�QUQUDE$���P(@$PA p ���/w�5�뮻����W�U���������][�׿ۯ�������/w�5�뮻����W�U���������][�׿ۯ��������/w�5�뮻����W�U���������][�׿ۯ�������Ј�*E�D(�(�*	Q"Q"DE$�� P) �QE p ���/w�պ�.���}�W�������ݻ��]\����k��������/w�պ�.���}�W�������ݻ��]\����k���������/w�պ�.���}�W�������ݻ��]\����k��������O�)D�OD
'Ǩ*N"�"D9$��P$�g�8� p ������ֻ�����8W������1ݻ���a]��?�q���������ֻ�����8W������1ݻ���a]��?�q����������ֻ�����8W������1ݻ���a]��?�q������                                   p �������������������������������������������������������������������������������������������������������������������������������                                   p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p ��������������������������������������������������������������������������������������������������������������������������������         �           �      p ������������������������������_��������������������������������������_���������������������������������������_�����������	   � @    @ �  �    H      �     p �����������������������������_�������������������������������������_��������������������������������������_�����������	   � @    @ �  �    H      �     p �����������������������������_�������������������������������������_��������������������������������������_�����������	��8�`g��`�����q�`k"��J���g<  p ���c1�}����Lq�mN4�>c�4㟔����}�_N3��������c1�}����Lq�mN4�>c�4㟔����}�_N3���������c1�}����Lq�mN4�>c�4㟔����}�_N3��������	"�D��H��A@��,��"
,��L���J��(H�  p ����n�}o�]�[��m5�}~���]o�]�]w���_5��]�������n�}o�]�[��m5�}~���]o�]�]w���_5��]��������n�}o�]�[��m5�}~���]o�]�]w���_5��]������	"�|�@H���@��肁>z�@H�"����(H�  p ����o�}��]�X0�Ut}~���A��A��w��U_u��]�������o�}��]�X0�Ut}~���A��A��w��U_u��]��������o�}��]�X0�Ut}~���A��A��w��U_u��]������	"�@� H��@���� �� H�"����(H�  p ����o�}߷]�[�Uu�}~�u�_߷_��w��U_u��]�������o�}߷]�[�Uu�}~�u�_߷_��w��U_u��]��������o�}߷]�[�Uu�}~�u�_߷_��w��U_u��]������	"�D��H��Q@D�(��"�(��H�����(H�  p ����n�}o�]�[���u�}~�u�]o�]�Yw���_u��]�������n�}o�]�[���u�}~�u�]o�]�Yw���_u��]��������n�}o�]�[���u�}~�u�]o�]�Yw���_u��]������	�8�`'�� D�ȂAyȜ`(������G<� p ����q�}����\p߻v7}��7c��c���~�_v;��������q�}����\p߻v7}��7c��c���~�_v;���������q�}����\p߻v7}��7c��c���~�_v;�������   �    �                �           p ��������������������������}��������������������������������������}���������������������������������������}���������������                       �           p ����������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p ���������������������������������������������������������������������������������������������������������������������������������������������������������������������� ��                                      ?����������������������������������������������������������������������������������������������������������������������������� ����������������������������������������������������������������������������������������������������������������������������������������������������������������������� �������������������������������������������                                       ��������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         ������������������������������������������������������������������������������������������������������������������������������