��`  ��#                                                                                                                                                                                                                                         ����������������������������������������������������������                                                                                                                                                                              ������������                                  ?�����������           ?�����������������������������������                                                                                                                               ����������������������������������������������������������                                                                                                                                                                              ����������������������������������������������������������                                                                                                        8                                                                     ����������������������������������������������������������                                                                                                        8                                                                     ����������������������������������������������������������                                                                                                        8                                                                                �����������������������������������           ������������                                  �����������                                              8                                                                     ����������������������������������������������������������                                                          ������������                                  ?�����������                                                          ����������������������������������������������������������                                                                                                        8                                                                     ����������������������������������������������������������                                                                                    ����������������� 8                                                                     ����������������������������������������������������������                                                                                                      8                                                                     ����������������������������������������������������������                   0                                                     0                      8                              0                                   ����������������������������������������������������������             1�   0  �                                               1�   0  �                      8                        1�   0  �                                   ����������������������������������������������������������             0    0  �                                               0    0  �                      8                        0    0  �                                   ����������������������������������������������������������             0|y�;||�|                                            0|y�;||�|                   8                        0|y�;||�|                                ����������������������������������������������������������             7�v́�v�6m�f                                            7�v́�v�6m�f                   8                        7�v́�v�6m�f                                ����������������������������������������������������������             1�f���f��m�f                                            1�f���f��m�f                   8                        1�f���f��m�f                                ��������������O�>fL�3�I�L���������������������������������                                                                      1�f���f��m�f                   8                                                                     ��������������L�2fL�3�I�L���������������������������������                                                                      3�f͙�f��m�f                   8                                                                     ��������������a��pd���̒`���������������������������������                                                                      �fy��f|3m�|                   8                                                                     ����������������������������������������������������������                                                                                 `                   8                                                                     ���������������������������������������������������������                                                                             �    `                   8                                                                     ����������������������������������������������������������                                                                                                      8                                                                     ����������������������������                �������������                           �����������������                                                           8                                                                     ����������������������������������������������������������                                                                                                        8                                                                     ����������������������������������������������������������                                                                                                        8                                                                     ����������������������������������������������������������                                                                                                        8                                                                     ����������������������������������������������������������                                                                                                        8                                                                                �����������������������������������           ������������                                  �����������                                              8                                                                     ����������������������������������������������������������                                                          ������������                                  ?�����������                                                          ����������������������������������������������������������                                                                                                        8                                                                     ����������������������������������������������������������                                                                     ?�����������������������������������                                                                     ����������������������������������������������������������                                                                     �����������������������������������                                                                     ����������������������������������������������������������                                                                     �����������������������������������                                                                     