�a  �U�n               �0     m�    ` 0                               �0     m�    ` 0                               �0     m�    ` 0                               �0     m�    ` 0                               �0   � ` ` 0                               �0   � ` ` 0                               �0   � ` ` 0                               �0   � ` ` 0                                0   � ` ` 0                                0   � ` ` 0                                0   � ` ` 0                                0   � ` ` 0                               3ǜ�m��sl�Ǐ3�                              3ǜ�m��sl�Ǐ3�                              3ǜ�m��sl�Ǐ3�                              3ǜ�m��sl�Ǐ3�                              ��l��m�n�cm��ٶl                              ��l��m�n�cm��ٶl                              ��l��m�n�cm��ٶl                              ��l��m�n�cm��ٶl                               ߷��m�l�cm���l                               ߷��m�l�cm���l                               ߷��m�l�cm���l                               ߷��m�l�cm���l                                                                                                                                   �6�3m�l�cm���l                                                                                                                                                                                    ٶl��3m�l�a͛ٶl                                                                                                                                                                                    �3ǌ��m���1���3��                                                                                                                                                                                             `  �                                                                                                                                                                                                  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �                ��               �                                                               �                ��               �             ` 0                              ` 0            ���              ���              ���            ��              ��               ��            �                 �              �                            @                            ���@             ����             ���@          ���              ���             ���              @             �                  @           ��              ��              ��           � �            � �             � �          ?����            ����             ?����          @��             ��             @��         � <              �            � <          ����            ?���?�           ����         �����            �����           �����         � <              �@           � <            �            �                 �         ����?�           �?����           ����?�        �����            �����           �����           ��           ��               ��         �   8               �            �   8         ?�����          �����~           ?�����        ������          ������           ������         �   8              �            �   8          ��            0 �� `            ��         |������          �������          |������        ������          ������           ������                       0    `�                      ����           @���@          ����       ������~          �������         ������~        �������          �������          �������           �          @                  �         ����`            ����            ����`       �������          �������         �������       �������          ?�������         �������             a          @                    a        �����        ��������        �����      ��������        �������{��       �������      ���������        ����������       ��������                            ���                      ����� �        �����@��        �����       ?����������      ����������       ?��������      ���������       ����������       ��������              �             B��                      �������        �����0�        �����       ���������      ���������       ��������      ?���������       ���������       ?��������      @      ��             1�       @             ���������       �������        �������      ��������{��      ���������       ��������x      ���������       ����������       ��������      �       � �                     �       �      �� ��E��      �� ��@       �� ��D     ����������      ����?����      ��������     ���� ����       ��� �����      ���� ���         �  @ �          �8             �  @       ��  ����       ��  ��@        ��  ��     ���� �����      ?��� ����      ���� ���     ���  ����       ?���  ����      ���  ���         �    �          �            �         ��   ��|�       ��  ���       ��   ��     ���  ���|�      ���  ?��p      ���  ���     ���   ���       ���  ����      ���   ���             �         @  0  �                   ��   �<�       �   ��@       ��   �     ���   ����      ���   ���      ���   ���    ���   ���       ���   ����      ���   ���       0   `  �             @         0   `      �    ��\�      ��    �$      �    ��@    ���   ����     ���    ���      ���   ���    ��    ���      ���    ���      ��    ���       �     �            �           �          �    ��,�      ��    �       �    ��     ?��    ����     ���    ?��      ?��    ���    ��    ���      ���    ���      ��    ���            �                                 ?�     ���       ��    �	        ?�     ���    ?��    ��t      ���    ��       ?��    ��p    ?��     ���      ���    ��p      ?��     ���             �                               �     �     ?�@       �     �        �     ?�@    ��     ��      ��     ��       ��     ��    ��     ?��      ��     ��       ��     ?��           @ @                            @ @     ��     �@       �     ��        ��     �@    ���     ��      ��     ���      ���     ��    ���     ��      ��     ���      ���     ��              @                                 @    ��     �$       �      ��@      ��     �$   ���     ��      ��      ���     ���     ��    ���     ��      ��      ���      ���     ��                                                  �      �       ?�      ?�       �      �   ��      ��      ��      ��     ��      ��   ��      ��      ��      ?��     ��      ��                          @                   �      �       ?�      �@      �      �   ��      ��      ?��      ��     ��      ��   ��      ��      ?��      ��     ��      ��                                                   �             @�      ��     �          ��       ��      ��      ��     ��       ��   ��       �      ��      ��     ��       �            �         @                      �     �       �       ��      �       �       �   ��       ?�      ��      �      ��       ?�   ��       �      ��      �      ��       �                                                     �               �                �            ��       �      ��        �      ��       �   ��               ��               ��                      �                �                �    �               �                �            ��              ��               ��            ��               ��               ��                                                            ?�               �                ?�            ��              ��               ��            ��              ��               ��                                                              ?�               �                ?�            ?��              ��               ?��            ��              ��               ��                                                              �               �                �            ?��              ��               ?��            ?��              ��               ?��                                                                               �                             �               ��               �             ?�               ��               ?�             @                                 @              @�               �               @�             �               ��               �             �               ��               �                                                                �                �                �             �               ��               �             �               ��               �                                                            �                �               �             ��               ��               ��             �               ��               �             �                                 �              ��               �               ��             ��               ��               ��             ��               ��               ��                                                             �                �               �             ��               ��               ��             ��               ��               ��                                                             �                ?�               �            ��               ��              ��             ��               ��               ��                                                           �               ?�              �            ��               ��              ��            ��               ��              ��                               @                             �                ?�               �            ��               ��              ��            ��               ��              ��                               @                             �                �               �            ��               ��              ��            ��               ��              ��                                                               �                �               �            ��               ��              ��            ��               ��              ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ? `              |�               l0                                                                                                                                                                  1�              ��               `0                                                                                                                                                                  1�              ��               `0                                                                                                                                                                  1�o�             ���?�            l��π                                                                                                                                                                ?n�             �홶ـ           �6n�                                                                                                                                                                0l�             �͙�߀           m�7��                                                                                                                                                                03l�             �͙��            m�6�                                                                                                                                                                03l�             �͙�ـ           m�6l�                                                                                                                                                                0l�             |͏6�            l����                                                                                                                                                                                                                                                               