�bb  (6dM             �      ��     � �                          �      ��     � �                          �      ��     � �                          �      ��     � �                          �      �      � �                          �      �      � �                          �      �      � �                          �      �      � �                                �      � �                                �      � �                                �      � �                                �      � �                          <q�<ݳ<�3<�<�8                         <q�<ݳ<�3<�<�8                         <q�<ݳ<�3<�<�8                         <q�<ݳ<�3<�<�8                         �f�0ٳfٳf�3fٰ                         �f�0ٳfٳf�3fٰ                         �f�0ٳfٳf�3fٰ                         �f�0ٳfٳf�3fٰ                         �fc�>ٞ~�~�0fٰ                         �fc�>ٞ~�~�0fٰ                         �fc�>ٞ~�~�0fٰ                         �fc�>ٞ~�~�0fٰ                                                                                                                   �f3 fٞ`�`�0fٰ                                                                                                                                                                ٳf�0fٌfٌf�3fٰ                                                                                                                                                                ��<q�>ٌ<�<�<�3l                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             �          ��          H     ��                      ��          H     ��          p           ��                                          ��                            ��         ���         $�     ���                     ���         $�     ���         p           ���                                         ���                           ����       ����       I     ����                    ����       I     ����        p           ����                                        ����                          �����      �����      �      �����                   �����      �      �����       p           �����                                       �����                          ������     ������             ������                  ������             ������                  ������                                      ������                         �������     ������            ������                  ������            ������                  ������                                      ������                         �������     ?������             ?������                  ?������             ?������                  ?������                                      ?������                         �������     ������             ������                  ������             ������                  ������                                      ������                         �������     ������             ������                  ������             ������                  ������                                      ������                         ������     ������           �������        �8        �������           ������          ������                                      ������             ����*��     ��_����     ¡S���             �������        �8        �������             ������     
��J����     ¡Q��                          @        ¡��                         ������     5 ��             �������        �8        ���c���             ����*��     UUEUUP     5 �t             UUQTUUU                                     UUUUUUT     �������     `����             �������                  ���             UUUUUUT     �������     `����             �������                    #�                           �������     �������            �������                  �������                        �������                         �������                                                  �������     �������             ������                  �������                         �������                         ������                                                  �������     ������             ������                  ������                         �������                         ������                                                  �������     ?������            ?������                  ?������                        �������                         ?������                                                  ������      ������            ������                  ������                        ������                          ������                                                   �����      �����       $�I$� ������                  �����       $�I$�              �����                          ������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             �          0         >`           �                                                                                                                                            �  �        �         c`           �                                                                                                                                            �  �        �         ``           �                                                                                                                                            ��|�        �Ǜ        `|�ǀ       �><                                                                                                                                          �v�        0l�        `v��l�       ٻf                                                                                                                                          ��f�        ��        `f��o�       ٳ~                                                                                                                                          ��f�        �l        `f��l        ٳ`                                                                                                                                          ��f�        �l�        cf��l�       ٳf                                                                                                                                          ��f`        3癀       >fǛg�       �3<                                               