��d  �	 
    ���������������������?������ � ���?��� � ���   � � ���   � � ?��   � � ����    � ������   ���                 
 ��� ( ��������� ( ��������� ( ��������� ( ��������� ( ���������)���������� ( ��������� ( ��������� ( ��������� ( ������                                                                                                                                                    C  ���������         ���������������������������         ����������������������������  |a� ����������������������������  �a� ���������������������������   �<s� ���������������������������3<�<s� �����������������������������f�f� ��������������������������� Ϟ~�f� ��������������������������� ٞ`�~m� ���������������������������ٌf��m� �����������������������������<~�a� ���������������������������         ���������������������������         ���������������������������         ������������������            C  ���������         ���������������������������         ���������������������������  >0߀���������������������������  c0� ���������������������������  `9� ����������������������������`9� �����������������������������o3?� ���������������������������ϳc3?� ���������������������������ٳc?6� ���������������������������ٳga�� ���������������������������珟?a�߀���������������������������         ���������������������������         ���������������������������         ������������������            C  ���������         ���������������������������         ���������������������������0 0  �   ���������������������������0 0  �   ���������������������������0 8  �   ���������������������������7�3�<������������������������������7m�3f͛�����������������������������6f33`͛3 ���������������������������6c33`͛1����������������������������6m�7f͛6����������������������������6g<l�3����������������������������         ���������������������������         ���������������������������         ������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        