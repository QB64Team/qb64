�/a  �W�f                    �       0`   �                                       �       0`   �                                       �       0`   �                                       �       0`   �                                      3 � `     0   �                                      3 � `     0   �                                      3 � `     0   �                                      3 � `     0   �                                      0 � `     0   �                                      0 � `     0   �                                      0 � `     0   �                                      0 � `     0   �                                      0<�p<x��l��m�                                      0<�p<x��l��m�                                      0<�p<x��l��m�                                      0<�p<x��l��m�                                      fٳ`�6lكlm�                                      fٳ`�6lكlm�                                      fٳ`�6lكlm�                                      fٳ`�6lكlm�                                      ~߰`>��6g���m�                                      ~߰`>��6g���m�                                      ~߰`>��6g���m�                                      ~߰`>��6g���m�                                                                                                                                                    `�0`f��6g� �m�                                                                                                                                                                                                           3fٳ`f͛6c�l9�                                                                                                                                                                                                           <�0>x��c�1�m�                                                                                                                                                                                                                        0                                                                                                                                                                                                                           �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 �                 �@                                ?��                 s�`                                ��                 ��                                0 `                 �                                ��                ��                               ��                ��                               ���                ���                               �                  ��            �                `x�                ����            �               ����               ����                               ��<                ��<                              �`                 ��8            (�               ���               ����            *�               ?�k��               s�����           �               ����               ����             �               0� �               ����           !���              �}�Ā             �����           ���              �����             �����@          -\�              ���߀             ���߀           \�              ��               ����          h �              `|� �@             ���� ��         ����             �������            �������         w�              �����             �����           �             �|  �              ��� ��        �  8             ��� ,�            '���� /�        &���             �����`            ��������        ��               ���� �            ���� �         �                `� @ �            ���� �        ��@&S.            ���&S*@           	����S+�        I��9��            ���9���           9�������        �x@&$            ����&#�           ����&'�           P$            �  P$@           ��� P#�       !�� fs7            ����fs7           ?���fs3�       i� y���           ����y���           ?���y���       -� &!            �����&!�           �����&!�        H   p!             �    p             ?��� p!�      �  ` 3�           ���` 3�           ���` 1�      �x  ���           ��������           ������      w�  �             ������ �           ����� �          @                 @             �� @ �     �  ��=�          a������=�          ���>��=�     &�  ����          ���������          ���>����     ��  � <�          ������ <�          ����� <|      �  � <�           `   � <�           �� >� <|     ��@  � >�          �?����� >�          ����>3� >�     I��  ����          I���������          I���>;����     �x@  � ~           ������� ~>          ������ ~>         � >               � >@          �� >#� >>    !��   ���`         !���������Q         !���|C���^    i�   � ~�         i������ ~�         i��|S� ~ހ   -�   ���@         -���������_         -��������     H    � >@          H    #� >`          H� |C� >^   �    �p?p        �������p?p        ���|g�p?�  �x    ��P        �x�������_        �x��|g��_�  w�    �w��        w�������w��        w������w��         �                �            � |G�    �     ���        � ���������       � �������  &�     � ?�       &� ������ ?߀      &� ����� ?�   ��     ��Ϡ        �� �������ϯ�       �� ���ϟ�Ͽ�  �     � �        �     O� �        � � ��� �  �@     �x�       �@ ������x�       �@ ���πx�� ��     ���       �� ���������      �� �������� �@     ?w��       �@ �����?w�߀      �@ � ?��?w�π �        �       �        �       �   ��  �� �      �8K�       �  �����8K�       �  ����8K�� �      �X��       �  ������X���      �  ���^�X��� �      W�W�       �  ����W�Wǀ      �  � ?��W�Wπ �       �       �      � �       �   � ǀ �      !8��0       �  ����!8��4@      �  ?���8��?� _      !D�4       _  ����!D�?�      _  ?���D�?� �      ����       �  ���������      �  � ������ _        �         _        �        _  > �  � � ?��     }�       ?�� ����}�@      ?�� ?���}�� ?��            ?�� �����      ?�� ?���� ?��     >����       ?�� ����>�����      ?�� � �>����� ?��               ?��               ?�� > �  � ?��     >q�       ?�� ����>q�       ?�� ��>q�� ~�     F       ~� ����F�      ~� ��F� ?��     <����       ?�� ����<�����      ?�� � ��<����� >�               >�              >� | �   � �      ��       �  ������       �  ������         ,p�           ����,p��          ���,p�� ��     =��]�       �� ����=��]��      �� ���=��]��          p                 p             � � p �       
���         ����
���         ���
���� ��      ��       ��  �������      ��  ������ |�     =��}�       |� ����=��}��      |� ���=��}��          �                 �            � � � �         ��L               ��N               ��K�       ��             ���            ��� ���     =��}�       ���     =��}��      ���     =��}��          �                  �                  � � ���     
���       ���     
���       ���     
���� ��`     ��       ��`     ���      ��`     ���   �     =��}�         �     =��}��        �     =��}��          �                  �                  � � ���     ��       ���     ��       ���     ��  ���     ,p�       ���     ,p�       ���     ,p�  p�     =��]�       p�     =��]�       p�     =��]�    �      p          �      p          �      p   ���     :q�       ���     :q�       ���     :q�  ��`     F       ��`     F       ��`     F    �     =����         �     =����         �     =����                                                      ���     �       ���     �       ���     �  ���            ���            ���             >����             >����             >����                                                       �      !=�        �      !=�8        �      !=�8  �      !E8       �      !E8       �      !E8  x��     ����       x��     ����       x��     ����                                                              ��{�               ��{�               ��{�  �      ����       �      ����       �      ����  |�     WW�       |�     WW�       |�     WW�           �                �                �          �p�               �p�               �p�  A�@     ���       A�@     ���       A�@     ���  >�     w��       >�     w��       >�     w��            �                 �                 �  ?��     ��`       ?��     ���       ?��     ���  ?��     � �       ?��     � �       ?��     � �  ?��     ���        ?��     ���       ?��     ���  ?��     �         ?��     � �       ?��     � �  �      �x?�       �      �x?`       �      �x?`  _      ��?�       _      ��?`       _      ��?`  �      �w�        �      �wߠ       �      �wߠ  _      �         _      �         _      �    �      �8��       �      �8��       �      �8��  �      �X�`       �      �X�`       �      �X�`  �      �?�       �      �?�       �      �?�  �      �>        �      �>        �      �>   �B     ��       �B     ��       �B     ��  ��     ��       ��     ��       ��     ��  �Z     ����       �Z     ����       �Z     ����  �      � |�       �      � ~�       �      � ~�   o��   ���         o��   ���         o��   ���    u�)    ����        u�)    ����        u�)    ����   �ր   ��         �ր   ��         �ր   ��    �     ��         �     ��         �     ��    [��    ��         [��    ��         [��    ��    �mJ@   ��         �mJ@   ��         �mJ@   ��     C���   ���          C���   ���          C���   ���     )     ��          )     ��          )     ��      ���  ?��           ���  ?��           ���  ?��     �[R�  ?��          �[R�  ?��          �[R�  ?��      ��h  ?��           ��h  ?��           ��h  ?��       J@   ?߀            J@   ?��            J@   ?��       5��B ��            5��B ��            5��B ��       {�Ԥ ��            {�Ԥ ��            {�Ԥ ��       ;�Z �            ;�Z ��            ;�Z ��        �  �             �  ��             �  ��        o��3�             o����             o����        ��)JR�             ��)M��             ��)M��        �ֵ�@             �ֳ�@             �ֳ�@         �   @              � �@              � �@         [���               [���               [���          �mj߀              �mj߀              �mj߀          C��r                C��r                C��r           )JR                )JR                )JR            ֵ�                 ֵ�                 ֵ�           �{�                �{�                �{�            �                  �                  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            0 �          � 0              ��     � 0                                                                                                                                                                           1�   0            l          �     ��      � 0                                                                                                                                                                           1�   0                      �     ��      � 0                                                                                                                                                                           1�<�><�          �7�}��> ��|�     �����<��>s���                                                                                                                                                                       1�f��݀         ��`͘6f �v�     ��6�����fm�`                                                                                                                                                                       1�~�3>ـ         ϶`͙�f ��f�     �����>��3fm��                                                                                                                                                                       1�`�3fـ         ٶ`͛6f ͛f�     ��6��f��3fm�                                                                                                                                                                        1�f��fـ         lٶ`ͻ6f ͛f�     ��6��f���fm�`                                                                                                                                                                       ><�3>ـ         �϶`|��>`��f`      �����>��3cͳ�                                                                                                                                                                        0                        ��             �                                                                                                                                                                                0                     �    �                                                                              