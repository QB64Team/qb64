�~]  X� 7                    �������������������                                      �������������������                                                        �������������������                                                        �������������������                                    0                   �������������������                                    0                   �������������������                                    0                   �������������������                                    0                   �������������������                                    0                   �������������������                                    0                   �������������������                                    0                   �������������������                                    0                   �������������������                                    0                   �������������������                                    0                   ������������������� p  B  >                            0                   ������������������� �  b  !   �                        0                   ������������������� �  b  !   �                        0                   ������������������� �9�RrH!g'�                        0                   ������������������� r R�H>H���                        0                   ������������������� 
= J�� H���                        0                   ������������������� 
E F�� H� �                        0                   ������������������� �E F� H���                        0                   ������������������� q=Bq G'@                        0                   �������������������                                    0                   �������������������                                    0                   �������������������                                    0                   �������������������                                    0                   �������������������                                    0                   �������������������                                    0                   �������������������                                    0                   ������������������� x                              0                   ������������������� �     �                       0                   ������������������� �  �   �                       0                   ������������������� ��s8�X�L���                    0                   ������������������� �"
D�eRR)$@                    0                   ������������������� �>z|QEUH�$�@                    0                   ������������������� � �@QEUD�%@                    0                   ������������������� �"�D!EH��%@                    0                   ������������������� yy8!D�%$��                    0                   �������������������                                   0                   �������������������                                   0                   �������������������                                    0                   �������������������                                    0                   �������������������                                    0                   �������������������                                    0                   �������������������                                    0                   �������������������                                    0                   �������������������                                    0                   �������������������                                    0                   �������������������                                    0                   �������������������                                    0                   �������������������                                    0                   �������������������                                    0                   �������������������                   �������������������                   ������������������                   ������������������                   ������������������                   ������������������                   