�i  $(� k 8                                              ?                       8                       G                       ;�                      �                      D                       ��                      |��                     ���                     �                       ���                     }�                     ���                     ��                      ���                     }�?�                    ����                    ��                     D���                    ;���                    |���                    G >                     ?��                    ���                   ?���                   8��                    z�?��                  ^����                   z�?��                  $�                    <���                   n���                  |����                   >�                   = >��                  / ?���                  = >��                   �                   ����                  7���~                  >����                  	  �                  � �                  � ���                 � ��                 	  �p                  @ ���                 � ���                 @ ���                 �                    @  �                 �  �>                 @  �                 �  ��                 �  ��                 �  ���                �  ���                @   p8                 �   q��                �   ��                �   q��                @                    �   ?�                �   �<                �   ?�                    ��                �   ��                �   �π               �   ���                    80                �    9��               x    ?��               �    9��                �                    �    ?�               x    �x               �    ?�                �    À                �    ��               �    ��               �    ��                H     0`                �     3�               �     ?�              �     3��               H                     z     �               �     ��               �     �               $     �                z     ��               �     �x               �     ��               $      a�               =      g�               o      �               }      g�                     `               =      �               o      �              }      ��                                   �     �              7�     ��              >�     �              	      �               �     ��              7�     �x              >�     ��              	       a�              @      g�              �      �              @      g�              �      `              @      �              �      �             @      ��             �                    �      �             �      ��             �      �             @      �              �      ��             �      �x             �      ��             @       a�             �       g�             �       �             �       g�                     `             �       �             �       �            �       ��                                 �       �            x       ��            �       �             �       �             �       ��            x       �x            �       ��             �        a�             �        g�            �        �            �        g�             H        `             �        �            �        �           �        ��            H                     z        �            �        ��            �        �            $        �             z        ��            �        �x            �        ��            $         a�            =         g�            o         �            }         g�                     `            =         �            o         �           }         ��                                �        �           7�        ��           >�        �           	         �            �        ��           7�        �x           >�        ��           	          a�           @         g�           �         �           @         g�           �         `           @         �   �       �         �  �       @         ��  p       �                    �         ���p       �         ��  p       �         ����       @         ���`       �         �� �       �         �_���       �         �����       @          a�  �       �          g� �       �          ���       �          g����                  @         �          � �       �          ���       �          ����                            �            �       x          ���       �          ?���        �           �          �           � �       x           ����       �           ���t        �                       �           ��r       �           ?��r�      �           ?���        H                       �           � ��      �           7� ��      �           >� w        H           	          z           � v        �           7� 7        �           >�         $           	          z           � 9�       �           7� ?�       �           >� p        $           	  0        =           � A�       o           7� ߠ       }           >�  @                  	           =           � `       o           7� `       }           >� 	�                  	  @       �          � �       7�          7� �       >�          >�         	           	          �          � `       7�          7� �       >�          >�         	           	          @          � `       �          7� 7�       @          >�         �          	           @          � �       �          7� �       @          >� p       �          	         �          � `       �          7� p       �          >� �       @          	          �          � �       �          7� �       �          >�         @          	          �          �        �          7� �       �          >�                    	           �          �  �       �          7� �       �          >�  �                  	   �       �          � �       x          7�  �       �          >�  `        �          	   @       �          �  �       x          7�  �       �          >� �        �          	   �        �          �        �          7� ~�      �          >�          H          	            �          �  9�      �          7�  y�      �          >�  '        H          	   !        z          �  t        �          7�  7�       �          >�          $          	           z          �  0        �          7�  ?        �          >�  p        $          	   0        =          �   �       o          7�  ��       }          >�  @                  	            =          �  �       o          7�  o�       }          >�                    	           �         �  @       7�         7�  �       >�         >�          	          	           �         �  @       7�         7�  �       >�         >�          	          	           @         �  �       �         7�  �       @         >�          �         	           @         �  �       �         7�  �       @         >�          �         	           �         �  �       �         7�  �       �         >�  �       @         	   �       �         �  �       �         7�  �       �         >�  �       @         	    �       �         �  �       �         7�  �       �         >�   �                 	    �       �         �  |       �         7�  G       �         >�   �                 	    D       �         �   �       x         7�  �       �         >�   �        �         	    �       �         �   �      x         7�   ��      �         >�   ��      �         	    �       �         �   � ��    �         7�   ����    �         >�   ����     H         	    �        �         �   {      �         7�   Ï�    �         >�   ����     H         	    @        z         �    >      �         7�   G�݀     �         >�   ���     $         	           z         �   �>      �         7�  �Հ     �         >�  ����     $         	    �      =          �  � >      o         ?� ��݀     }         ?� �� ��                  ��      =            �       o         ?�����     }         ?��� ��                 ���       �         � �       7�        �������     >�        q��� �      	           ��� ��     �        � �       7�        �����       >�        ��� �       	          ���         @        ?� �         �        �����         @        �p �         �         ��          `        ?��          �        ����          `        �`�          �        �           �        ?��           �       ���           �        �o�           @                    �                    �       ��            �       ��                                  ��  �              ?����������            �������q�             �       �             ������              �       ��            ���������?�             ?�������               �  �  �              ����������               �  �  �              ���������                       �              �������               �  � �              ������`              ��������               ������               ��������                                       �  �                  �  �                                                                 �                                              �                                              �    0                 �����                 �                                             ������                                        ������                                         �    <                                        �    4                                                                                                                                