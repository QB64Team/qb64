�l  �z��                 `                                              `                                              `                                              `                                             �` 0                                           �` 0                                           �` 0                                           �` 0                                            ` 0                                            ` 0                                            ` 0                                            ` 0                                           g�8<��ny����<��<                               g�8<��ny����<��<                               g�8<��ny����<��<                               g�8<��ny����<��<                               3lٰf��l��m���f                               3lٰf��l��m���f                               3lٰf��l��m���f                               3lٰf��l��m���f                               �o�0f�������0>͛~                               �o�0f�������0>͛~                               �o�0f�������0>͛~                               �o�0f�������0>͛~                                                                                                                                       �l03f�����͛0f͛`                                                                                                                                                                                           �lٰ3f́�l͛m�0f͛f                                                                                                                                                                                           g�<���fy���0>��<�                                                                                                                                                                                                                                                                                                                                                                                                                           �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ?��                ��                ��                                                                                                                                                                       � |                �               | �                                                                                                                                                                      x  �             �                �  <                                                                                                                                                                     �   8                 �             8   �                                                                                                                                                                                     0                 �    `                                                                                                                                                                    0    �            �                                                                                                                                                                                         �     `                �                                                                                                                                                                                                          `           0     �                                                                                                                                                                                   0                 �      `                                                                                                                                                                                   @                                                                                                                                                                                                 �          �                                                                                                                                                                                         �       `                �                                                                                                                                                                                                          @                                                                                                                                                                                                                             �                                                                                                                                                                                                  @        @                                                                                                                                                                                                   �                                                                                                                                                                                          @                                                                                                                                                                                                   �        �                                                                                                                                                                                         @         @                                                                                                                                                                                                 �                           �                                                                                                                                                                                                          @                                                                                                                                                                                                                             �                                                                                                                                                                                                           �                                                                                                                                                                                              @          @                                                                                                                                   @                                                           �                                                                                           @                                                  �                                         @                                                                                                           �                                                  �                                         @                                                                                                           �                                                                                      �      �                                                                                                                                                                                                �      �                                                                                                                                                                                    @           @                                                                                                                                                                                     @     @           @                                                                                                                                   @                                                 �     �                             �                                                                                                                  �                                                       �                             �                                                                                                                                                                                                      @                                                                                                                               @                                                                       @                                                                             @                                                  @                                                                                          �                                                            @                                                  �                  @                                                                       �                                                            �                  @                               �                  �                                                                        �                                                            �                  �                                                  �                  @                                       @            @                                                                              �                  @                                                 �                                       @            @                                                                                                �                                                                                        @            @                                                                                                                                                                                        @            @                                                                                                                                                                                         �                                                                                                                                                                                         �          �                                       @                                                                                                   �                  �            P                �          �      �             0                 �                  @                               �                               P                 �                 `            T                �          �     `             8                 �                  �                               �                  `             �                 �                 �            �                �          �     �             t                 �                 �                               �                  �             �                 R                 �            �          @                    �            t                 �                 �                                                 �            D                 �                 �           T          @     �               �            �                 8                 �             @                                   �            D                 �                 @           T          @     $               `            �                 �                 �             @                                                �                 H                 .�           �          @     ,H               .�           ��                �                 <             �                                                ��                .                 ]<           ��         @     /               ]�           �>                ��                >C�            �                                                �                ^��                ��          _�         @     \��              ��          ���               ;o�               |�           �                                 8|            ��               5?��              t��          _��        @     �?��            v��          �>               ~��<               ���           >                0 �                p�           
'��               �_��              ���         
���        @     ���            ����         @��              s���             �            �               0 �               �            
8?��             z ���             Ӄ��         
����       @    r���           ����         @               � <<             �  ��                          `  <              �  �          W���              ����             �|��        w���       @    �����           ����        �  ��            �  À            �              �              �  �             �            `~��            ��?��            N���        p���      @    ������          o���        �              �   <p            �   ��                         �   <                �         (����            ����            ����       *����      @    �����          ߀���           �           �   �            (   8            �            �   �                        (� ��           S� <?�            @ ���       *� ���     @    � ?��          �� ���       @   p           �    q�           T   �        @                   p               �        Q�  ���           �� ���           @ �       U�  ���     @    �� ���         � ��       :@   �           9    8           �    8�       @   �                               8        z  �           ��  <�            �  ���      ~  ��     @    %�  ?��         �  ���      �    q�          ڀ   �           
                p            �   �                        z   ���           I�  ��           @�  ?�      ~   ���          I�  ��     �     �  ��            0           ��    8�                �                         �    8           @     �       =   �          �   q��          ��  ��       ?   ��           P�   ��     �     �  ��        P    �           @    0                �          �           @               �             =   ��           �   ?�          �   8��      ?   ��            �   ��     �     �   ?��       P     0           @     �                             0           @     �                       �   q�           z   ��          �   �      �   �            ~   ��     �     �   ��       (                 �     0           �     �                             0           �     �      @�   <           z    8�          �    ��      �   �            ~    ?�     �     �    ��       (                  �                 �            @                                   �            @@   �           =                �    �      �   �           ?    �     @      �    �                         P                 @            @                                  @            �@    0           =     �           �           �    <           ?     �     @      �    �                         P                 @            �                                  @            ��               �                 z     �      �               �    0     @      ~     �       
                  (                  �            �                                                �                 �              @  z            �               �         @      ~     @       
                  (                  �                                             @               �                 @              �  =            �               �                 ?     �                                           P                                             �              �               @ @                =            �               �                 ?     �                                           P                            @                              �               � �                �           �               �                 �    �       �                 
                  (             �               �                              �               � �                �           �               �    @           �           �                 
                  (             �               �                               �                �                @            �               �    @           �           @                                                @                                              �                �                @      �      �                �    �           �           @                                                @                                              z                �                 �      �      ~                �    �           �            �                 �                 
                               �                              z                �             @   �      @      ~    @           �               �            �                 �                 
                               �             @                =                 �             �   �      @      ?    @            �               �            P                 @                                               @             �                 =                 �                �             ?    �      �      �               �            P                 @                                                @                              �                z                �             �   �      �      ~               �            (                  �                 �                                                �          @  �                 z                �            �         @      ~               �            (                  �                 �          @                                      �          @  @                 =                 �            �         @      ?                �                              P                 @          @                                     @          �  @             @   =                 �            �                ?          �      �                               P                 @          �                @                    @          �  �             �   �                 z            �               �         @      ~   @         
                  (                  �          �                �                                  �             �   �           @     z            �               �                 ~   �         
                  (                  �                          �               @                  �                @           �     =            �               �                 ?   �                                             P                                         �                 �                @                =            �               �  @             ?                                                P                                                          �                �                �      �     �                �  �             �           �                 
                  (             �                                             �                �                 �      @     �  @             �               �           �                 
                  (             �                                               �                �                 @             �  �        �     �               �           @                                                @                                               �                �                 @            �          @     �               �           @                                                @                                               z                �                 �            ~                �          �     �             �                 �                 
                               �                              z                 �                 �            ~               �          @     � @           �                 �                 
                                �                              =                  �                 �            ?                �                 � �           P                 @                                                @                               =            @     �                 �            ?                � @              �            P                 @                                           @     @                               �           �     z                 �       �     �`               ~�              �            (                  �                 �                         �                        �        @    �                 z                 �             ��          �     ~               �            (                  �                 �        @                                         �        @    @                 =                  �            �           @     ?                �                              P                 @        @                                        @        �    @                 =                  �            �           0     ?           �     �`                              P                 @        �                                        @        �    �                 �                 z            �                �           0     �            
                  (                  �        �                                                      �                                   x        �    �                �                ~             
                  (                  �                                                                                                            0    �            �                     8                                                 @                                                                                                                                 0                 �    `                                                                                                                                                                    �   8                 �             8   �                                                                                                                                                                     x  �             �                �  <                                                                                                                                                                      � |                �               | �                                                                                                                                                                       ?��                ��                ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      � `�  ��         ̀`             �         0                                                                                                                                                              0    ��         l `�             0     0                                                                                                                                                                 0    ��          `�             0     0                                                                                                                                                                 1�n�><��;`<��<     �|�y�<��y�      ��͹��3π                                                                                                                                                            1��lٻ�����f     ͳv�Ͷf���      ͳ3m�m�7m�n�                                                                                                                                                            1��lٳ>����>͛~      m�f���~��͘      3?m��3�f6l�                                                                                                                                                            1��lٳf����f͛`      m�f���`�f͘      30m�3c6l�                                                                                                                                                            1��lٳf���`f͛f     m�f�ͶfͶ͘      �3m�m�6m�l�                                                                                                                                                            1��f�3>��30>��<     ͟f`y�<��y�      �m�͙�g3��                                                                                                                                                                                                                                                                                                                                                                                      �        >                                                                                 