��b   ��M                                                                            �������������������                            �������������������                                                                            �������������������                                                                                                                        �������������������                            �������������������                                                                                                                          �������������������                            ?�������������������                            @                                              @                                              ?�������������������                            |                                              ��������������������                            ��������������������                            |                                              �                                             �������������������                           �������������������                            �                                             �                                             �������������������                           �������������������                           �                                             �                                             �������������������                           �������������������                           �                                             �                                             #�������������������                           #�������������������                           �                                             �                                             C�������������������                           C�������������������                           �                                             x                                              ��������������������                            �                                             {����   ���   ����                           >�                                             A�������������������                           A                                             >�m��rI$�6�m�$�I#m��n                           }�                                             ��������������������                           �                                             }�����   ���   ����                           ��                                            ?�������������������                                                                        ������   ���   ����                          ��                                            �������������������                          @                                            ��m��rI$�6�m�$�I#m��n                          �                                             ��������������������                          �                                            �����   ���   ����                          �                                             !��������������������                          !                                             �����   ���   ����                          �                                             C��������������������                          B                                             �#m��rI$�6�m�$�I#m��n                          x                                              ���������������������                           �                                             x����   ���   ����                          >�                                             A��������������������                          A                                             >�����   ���   ����                          }�                                             ���������������������                          �                                             }�#m��rI$�6�m�$�I#m��n                      �� ��                                         ��?��������������������                                                                   �� ������   ���   ����                      ����                                          l��������������������                       ��@                                         ��������   ���   ����                      ����                                          ������������������������                      ���                                         ����I#m��rI$�6�m�$�I#m��n                     ����                                         ���(!���������������������                      ��!                                         ���� ����   ���   ����                     �{￼                                         ^@�C���������������������                     �{�B                                         �{￼ ����   ���   ����                     �{�x                                         � d����������������������                     �{�x�                                         �{�zI#m��rI$�6�m�$�I#m��n                     s�{�}�                                         w{�u���������������������                     � _x                                         w�{�}� ����   ���   ����                     ��{���                                         �o{������������������������                     7� �                                         ��{��� ����   ���   ����                    �����                                        ��������������������������                     z  �                                         �����I#m��rI$�6�m�$�I#m��n                    ������                                        A����?���������������������                     �   w�                                        ������ ����   ���   ����                    =�{��                                        ��{�����������������������                    �   /�                                        ��{�� ����   ���   ����                    ���x                                        �����������������������                    � {�/`                                        ����}�ܒI$���m�$�H�m�ܒI$�                    ��C��                                        ��C؏���������������������                    `{��                                        �������   ����  ����                       =�H����                                        2H���o���������������������                    �7 z�                                        ?�������   ����  ����                       ;�L ��                                        $�L x�/���������������������                     � g�                                        ?�� ��ܒI$���m�$�H�m�ܒI$�                    w�0 ?�                                        i�0 �?���������������������                    � ���                                        �� ����   ����  ����                       ��@ �                                        ��@�����������������������                    ���@                                        ��� ����   ����  ����                       ������                                        ���?�����������������������                    4 ?p                                         �������ܒI$���m�$�H�m�ܒI$�                   �� �'�                                       �� �����������������������                    x �                                        �� �?���   ����  ����                      �� �                                        '� ?#����������������������                    � ?                                        �� ����   ����  ����                      � �                    >                    O ^ ����������������������                    �0 ^                   >                    �8 �m�ܒI$���m�$�H�m�ܒ$�                   �� @                    Y                    �  ��������������������>�                   �@  �                    ��                   �� @���   ����  ���� ��                   �� >�                    �                   � A8�������������������A?�                   �p A8                   ��                   �� >����   ����  ������                    }�                   ��                    �p������������������� ��                     � �p                   ��                   � }�[m�ܒI$���m�$�H�m�ܓ��                   � ��                   @�                   �c��������������������@_�                   �``                   ��                   �� ������   ����  ������                   ���                    �`                   �����������������������_�                   � �                   A�                   �������   ����  ������                   � �                    ��                    ������������������������                   ���                    `                   ����m�ܒI$���m�$�H�m�ܓ��                    ��                    ��                    �!������������������������                      !                     `                    ������   ����  ������                   � �                    ��                   < C�����������������������                   ��B                     �                   �������   ����  ������                                            ��          ����������������������������������?�          �������������                    ��                       H�m�ܒI$���m�$�H�m�ܓ��          �������������                     c�                      /����������������������?�                      (                    ��          �����������������   ����  ������          �������������                     ?                       ?���������������������@�                      0                     ��          �����������������   ����  ���� ��          �������������                                            ?������������������������                                            >           �������������H�m�ܒI$���m�$�H�m�ܒ$�                     �                                 ������������?������������������������          ������������                                             �����   ����  ����                        �                                 ������������?������������������������          ������������                                             �����   ����  ����                        �                                 ������������?������������������������          ������������                                             �H�m�ܒI$���m�$�H�m�ܒI$�                     �                                 ������������?������������������������          ������������                                             �����   ����  ����                        �                                 ������������?������������������������          ������������                                             �����   ����  ����                        �                                 ������������?������������������������          ������������                                             �H�m�ܒI$���m�$�H�m�ܒI$�                     �                                 ������������?������������������������          �                                            $�6�m�$�I#m������   ����  ����                        �                                 ������������?������������������������          �                                              ���   �������   ����  ����                        �                                 ������������?������������������������          �                                              ���   ��ͷ$�I#m��rI$�6�m�$�I#m��n                     �                                 ������������?������������������������          �                                            $�6�m�$�I#m���   ����   ���   ����                     �                                 ������������?������������������������          �                                              ���   ����   ����   ���   ����                     �                                 ������������?������������������������          �                                              ���   ��ͷ$�I#m��rI$�6�m�$�I#m��n                     �                                 ������������?������������������������          �                                            $�6�m�$�I#m���   ����   ���   ����                     �                                 ������������?������������������������          �                                              ���   ����   ����   ���   ����                     �                                 ������������?������������������������          �                                              ���   ��ͷ$�I#m��rI$�6�m�$�I#m��n                     �                                 ������������?������������������������          �                                            $�6�m�$�I#m���   ����   ���   ����                     �                                 ������������?������������������������          �                                              ���   ����   ����   ���   ����                     �                                 ������������?������������������������          �                                              ���   ��ͷ$�I#m��rI$�6�m�$�I#m��n                     �                                 ������������?������������������������          �                                            $�6�m�$�I#m���   ����   ���   ����                     �                                 ������������?������������������������          �                                              ���   ����   ����   ���   ����                     �                                 ������������?������������������������          �                                              ���   ��ͷ$�I#m��rI$�6�m�$�I#m��n                     �                                 ������������?������������������������          �                                            $�6�m�$�I#m���   ����   ���   ����                     �                                 ������������?������������������������          �                                              ���   ����   ����   ���   ����                     �                                 ������������?������������������������          �                                              ���   ��ͷ$�I#m��rI$�6�m�$�I#m��n                     �                                 ������������?������������������������          �                                            $�6�m�$�I#m���   ����   ���   ����                     �                                 ������������?������������������������          �                                              ���   ����   ����   ���   ����                     �                                 ������������?������������������������          �                                              ���   ��ͷ$�I#m��rI$�6�m�$�I#m��n                     �                                 ������������?������������������������          �                                            $�6�m�$�I#m���   ����   ���   ����                     �                                 ������������?������������������������          �                                              ���   ����   ����   ���   ����                     �                                 ������������?������������������������          �                                              ���   ��ͷ$�I#m��rI$�6�m�$�I#m��n                     �                                 ������������?������������������������          �                                            $�6�m�$�I#m���   ����   ���   ����                     �                                 ������������?������������������������          �                                              ���   ����   ����   ���   ����                     �                                 ������������?������������������������          �                    ��������������            ���   ��ͷ$�I#m��r@                                  �         ��������������          ������������?����������                       �                                            [m�$�H�m�ܒI��   ������������������                     �         ?��������������          ������������?����������                       � ��  ��           @                       ��  ��   ��   ����?��������������            �   �� �         ��������������          ��� ���� ��?����������                       � � �              �                       �� ���� ͷ$�I#m��r��������������            ��   �� �         �                        ��  ���� ��?�����������������������          �  �             ��������������          [l��H�m���I��   �����                         ��   �� �        �                        ��  ����  ��?�����������������������          �  �    �         ��������������          ��� ���� ��   �����                         �      ��        �                        ����������?�����������������������          ���  ��@         ��������������          ��  �� ��H�m�ܒI$��                         �      ��        �                        ��/�������?�?���������'��������������          �/��  ��          '��������������          [g� H�l �I�����   �                         �      ��        �                        ��O��������?���������G��������������          �O��  ��         G��������������          �  �� ������   �                         p      ��        p                        �����������?����������                        � ���  ��          �                        �p  �� ��H�m�ܒI$�p                         >�       ��        >�                        ����������?���������                        �A��  ��         A                        [>� H�l  �I�����   >�                         }�       |�        }�                        �����������?���������                         ��      �         �                         }�  ����|�����   }�                         ��       >�        ��                        �?���������?��������@                        �       �        @                        ~��  ����>�H�m�ܒI$��                        ��       �       �                         ����������?���������                        �@      ��        �                        Y��$�H�m��I�����  �                         �        ��       �                         ����������~?��������                         ��      �B                                 {�   ����������  �                         �        ��       �                         �!���������>?��������"                         �!        �"        "                         wހ  ������H�m�ܒI'�                         �        ��       �                         �C���������?��������D                         �B        |        D                         O��$�H�m�܃������  �                         x        ��       p                         �����������?���������                         ��        >
         �                         _{�  ����������  p                         >�         ��       >�                         ������������������                         �               A                         >��  ���� ��H�m�ܒI>�                         }�         }�       }�                         �������������������                          �        �       �                          }��$�H�m�ܐ}�����  }�                         ��         >�       ��                         !?�����������������@                         !         �      @                         �߀  ���� >�����  ��                         =��         |      �                          B�������������������                         B@        ��      �                         =���  ���� |H�m�ܒI�                          {�          �      �                          ������������A�������                          ��        �A                                {�m�$�H�m�ܒ����� �                          ��          �      �                         !����������� �������"                         !          � �     "                          ����  ���� ����� �                         �          �     �                         C�����������������D                         B          |@     D                         ���  ���� ��m�ܒO�                         �x          ��     p                          ������������?�������                          �          >       �                         �{m�$�H�m�ܒA������ p                         ��           ��     >�                         A�����������������                         A               A                         ����  ����  ������ >�                         }�           }�     }�                         �������������������                          �          �     �                          }���  ����  }��m�ܒ}�                         ��           >�     ��                         !?�����������������@                         !           �    @                         ��m�$�H�m�ܒH>����� ��                         =��           |    �                          B�������������������                         B@          ��    �                         =����  ����  }�����                          {�            �    �                          ��������������A�����                          ��          �A                              {���  ����  ��m�ܓ�                          ��            �    �                         !������������� �����"                         !            � �   "                          ��$�6�m�$�I#m������                         �            �   �                         C�����������������D                         B            |@   D                         �  ���   ��������                         �x            ��   p                          ��������������?�����                          �            >     �                         �x  ���   �����m�ܟp                         ��             ��   >�                         A�����������������                         A               A                         ��$�6�m�$�I#m�������>�                         }�             }�   }�                         �������������������                          �            �   �                          }�  ���   ���}����}�                         ��             >�   ��                         !?�����������������@                         !             �  @                         ��  ���   ���>��I"��                         =��             |  �                          B�������������������                         B@            ��  �                         =��$�6�m�$�I#m��|  �                          {�              �  �                          ����������������A���                          ��            �A                            {�   ���   ����  �                          ��              �  �                         !��������������� ���"                         !              � � "                          ��   ���   ����I'�                         �             � �                         C�����������������D                         B              |@ D                         �I$�6�m�$�I?m��� �                         �x           �  �� p                          ����������������?���                          �              >   �                         �x   ���    ������ p                         ��          @@   �� >�                         A����������������                         A               A                         ��   ���   @�����I>�                         }�          �    }� }�                         ������������?������                          �              � �                          }�I$�6�m�$�I�-��p}� }�                         ��             >� ��                         	?���������� �����@                         	               �@                         ��   ���   ���>� ��                         ��              ��                          	���������� ������                         	@             ��                         ��   ���   ����I�                          �               ��                          	����������� �����                          	�             �                          �rI$�6�m�$�I ��r��                          �               ��                          	����������� �����"                          	               �"                          ��   ���   �����                          �               ��                          	����������� �����D                          	               qD                          ��   ���   ����O�                          �                �p                          	����������� ?������                          	           �    1 �                          �rI$�6�m�$�I�-��rN�p                          �            @   �>�                          	�����������������                          	           @    A                          ��   ���   @����>�                          �            �   �}�                          	������������������                           	                �                           ��   ���    �����}�                          �               ���                          	�����������������@                          	               @                          �rI$�6�m�$�I?m��rN���                          �                ��                           	������������������                          	                �                          ��   ���   ������                           �                ��                           	�����������������                           	                                           ��   ���   ������                           �                ��                           	�����������������"                           	                "                           �rI$�6�m�$�I#m��rN��                           �                �                           	�����������������D                           	                D                           ��   ���   �����                           �                �p                           	������������������                           	                �                           ��   ���   �����p                           �                ��                           	�����������������                           	                                           �rI$�6�m�$�I#m��rN��                           �                ��                           	�����������������                            	                                            ��   ���   ������                           �                �                           	�����������������@                           	                @                           ��   ���   �����                           �                �                            	������������������                           	                �                           䍶�m�$�H�m�ܒI$���                            �                �                            	�����������������                            	                                            �����  ����   ��                            �                �                            	�����������������                            	                                            �����  ����   ��                            �                �          8                 	�����������������                            	                          8                 䍶�m�$�H�m�ܒI$���                            �                �          |                 	�����������������                            	                          |                 �����  ����   ��                            �                �          �                 	�����������������       �                  	                          �                 �����  ����   ��       �                  �                �          �                 	�����������������       � (�                	                          �                 䍶�m�$�H�m�ܒI$���       � 8�                �                �      �  �                 	�����������������       ��                	                      �  �                 �����  ����   ��       ��                �                �      �  �                 	�����������������       ��                	                      �  �                 �����  ����   ��       ��                �       �       �      ?�  ~                 	�����������������       ��                	                      ?�  ~                 䍶�m�$�O�m�ܒI$���       ��                �               �      � 8                 	��������?��������       �C�                	                      � 8                 �����  ?���   ��       �C�                �              �      �                   	����������������      ���                	                      ~�                   �����  ���   ��      ���                �               �      �  �               	����������������      ��	�                	                      x�  �               䍶�m�$�`m�ܒI$���      ��	�                �       @       �      ��x���               	����������������       �
�                	                      ��x���               �����  @���   ��      ���                �               �      �y���               	����������������       �
?�                	       @              �y���               �����  @���   ��       ����                �               �      ?�`
��               	����������������      @�?�               	       @              ?�`��               䍶�m�$�@m�ܒI$���      @���               �               �      �  �               	����������������      ��?�@               	       @              �   |               �����  @���   ��      �?�?��               �               �      �  �               	����������������     ��	�                	       @              �   <               �����  @���   ��     ����               �               �       p  �               	����������������     	����              	                       p  <               䍶�m�$�`m�ܒI$���     	�����              �               �       � ��               	����������������     ����                	                      �  �               �����  ���   ��     ���"                �                �        � ��               	��������?��������     ��&r�                	                       �  �               �����  ?���   ��     ��r                �       �       �        � ��               	�����������������    ��g*?�                	                       �  G�               䍶�m�$�O�m�ܒI$���    ��g*<@                �                �        p ��               	�����������������    ��7�$o�                	                        p  ��               �����  ����   ��    ��7�&l�               �                �     8 � �               	�����������������     �?�gO��               	                     8     @               �����  ����   ��     �<~gNF�               �                �     | �   <               �����������������     ��G��                                    |      <               䍶�m�$�H�m�ܒI$���     �>G��               �                �     | �                  9�����������������     ��F�3�               9                     l                    �����  ����   ��     �F�3�               �                �     �8�  ǀ              y�����������������     ������                y                     � �  ǀ              �����  ����   ��     ��ҟ����              �                �     �|�  �              ������������������     ���t��                �                     �    �              䍶�m�$�H�m�ܒI$���     ���t���              �                �    �|�  �              ������������������     ����	O�             �                    �    �               �����  ����   ��    ��?�	O�              �                �      |�  ��             ������������������    ������ `             �                           p�              �����  ����   ��    �������              �                �    �8    ��             ������������������     �����L              �                    �     ��              �rI$�6�m�$�I#m��rN�    ������L�              �                �         �p             ������������������     �����              �                          �p              ��   ���   �����    �����p              �                �         �p             ������������������     �����?�             �                          �p              ��   ���   �����    �����?�             �                �          8             /������������������     ��������             /�                          8             �rI$�6�m�$�I#m��rN�    ����d����             0�                �         8             O������������������     ���`��              O�                          8             0��   ���   �����    �{�` ��8             p�                �      �?�               �������������������     �_D�?�              ��                      �?�               p��   ���   �����    �D�?�             ��                �     �?� p            ������������������     ��J�              �                       ?�               ��rI$�6�m�$�I#m��rN�    �J�             ��                �     �?� �             ������������������     ��D���             �                     ?�               ���   ���   �����    �D��            ��                �    <� �             ������������������     ��`���             �                    < @                ���   ���   �����    <�G`�#�            ��   �           �      � �             /������������������    ��p?����            /�                       �  p             �v�rI$���m�$�I#m��rN�    ���p?�s��            ��              �    8 �  �             O�����������������    ���r�a���            O	                    8 H                 ����  ���   �����    ��Gr��#��            p�              �    8 �   �              ������������������    �?��3�����             �	                    8                    p���  ���   �����    �?�3����            >��              �    8  �  p             A�����������������    =�_#���            A	                !    8  �                 >���rI$��m�$�I#m��r^�   8=�#���            }��              >�    x    ��             ������������������    @!�"p�	            �	                A    8     ��             }����  ���   ����>�    x!�"qp�            ��|               }�    x   ��            ������������������    @�� �           �               �    8   ��             ���}�  ���   ����}�    x�� �           ���               ��    x    ��            ?�A���������������0    @���@��            A              0    8    ��            ����rI$��m�$�I#m��r��    x���@��           ��              ��    x p  �            � ���������������P    @���� a           @ �             P    8    �            ���`  ���   ������    x���� o           � �             �`    �  �  �� �           �����������������    �;����� !�           �@             �    8     ��            �6��  ���   �����`    �;���� /�          �  ��             ��    � �  �� �          A��?��������������!    �_���� ��          A               !    <     ��            ����I$��m�$�I#m��w��    �_�S����          |  {�             ��    � � �� �           ������������������B    �����@`�           � �             B         ��            |�{�  ���   �����    ��#��@`�          >�  =�             {�    � ��> �� �          A������������������    ����  0�          A �              �     �   ��            >�6�=�  ���   ����{�    �S�� 0�          }�  �   p          >��    ���>�� �          ������������������     �������          � �  �          A     �  ��            }���I$���m�$�I#m��>��    ������          ��  |              }�    ��p>� 9�         �������������������@    �G�7O��          ��              �@    �  � >           ���|   ���   ���}�    �G�H�?�         ��  �              ��     �� ?� 9�         ?���A�������������� �    ��� �            �A              �    �  ?� >          ��6��   ���   �����     ���	 ?�         �  �             ��     � �   � q�         ��� ��������������A     ��� �         @  | �            A      �   � ~          ����I$�6�m�$�I#m����     ��� �         �   �            �|     �     � q�          ������������������     ���0�          �  >@            �          � ~          � ���  ���   ����|     ���0�         �    ��            ��     ��       �         A����?�������������!     ����� �         A                !     �       �          ��6� ��  ���   �����     ������ ��         |    {�            ��     ��       �          �������������������B	     ����� �          �   �            B	     �       �          | ��{�$�6�m�$�I#m�Ͻ�     ������ ��         >�    =�            {�     ��     À         A�������������������     ��r� �         A   �             �     �      �          >� ��=�  ���   ���{�     ���r���         }�    �            >��     ��      ��         �������������������!     ��?
� �         �   �            A!      �      �          }��6� �  ���   �����     ���?
���         ��    |            }�     �  �   �         �������������������A     ��             ��            �A      �  �   �          �� ��|�m�$�H�m�ܒI}�     ����         ��    �            ��~     � �            ?�����A������������ �     � H�               �A            �      x �   �         �� ������  ����  ��~     � J��         �    �           ���     � �   <         ����| ������������A     � M�          @    | �          A       �   ?�         裸6�@���  ���� ���     � M�?�         �     �          �}�     � �   |          �����>������������     � BM�            �    >@          �       �   �         �  ���m�$�H�m�ܒK�}�     � BM� �         �      ��          ���     ?���   �         A�����?�����������!     ?�  �           A                !      ��   ��         �  �� ����  ���� ���     ?�� � ��         |      {�          ���     ?���  �          ������������������B     ?�              �     �          B      ��  ��         |�m�$� {���  ���� ���     ?�� ��         >�      =�          {��     ?�� �  �         A������������������     ?�  B           A     �           �      � �  ��         >����   =�m�$�H�m�ܒ_{��     ?�� B��         }�      �          >���     �|              ������������������      �  �           �     �          A       �    ��         }����   ���  ���� >���     �� ���         ��      |          }��     �>    > <        ������������������@     �     <             ��          �@      �    ?��         ���m�$� }��  ���� }��     ��  ?��        ��      >          ���     ��   � <        ?������������������ �     �      <               ��          �      ��   ���        �����   >m�$�H�m�ܒ���     ���  ���        �               ����     ��  � x        ������x�����������!      �       x        @      x��        !        ��  ���        ����   �  ��������     ���  ���        �       �        ����     ���  ��x         �������8����������"      ��    �x         �      8�@        "        ?�  �?�        �6�m�$�@��  ��������     ���  ���        �       �        ����     ���� �        A��������?���������.$      ��     �        A       �         .$        �����         �����   ��$�H�m�ܗ����     ��������        |       �        ����     �����> �         ������������������N(       ��    > �         �       �        N(         A������         }����   �  ��������     ���������        >�       �        q���     �ǃ�����        A������������������0 @     �ǀ   ��        A       �         �0 @       8����         >���m�$�H��  ����q���     ���������        }�        �        >���      ���  ��        ������������������  �     ���  ��        �       �        A  �       ���?�         }�����   @��$�H�m�ܾ���      ���������        ��        |        }���      ���� �       ������������������>       ���� �              ��        �"         �?� ��         ������  `}�  ����}���      ���������       ��        >        ����      ����� �       ?������������������~       ����� �               ��       B         �  ��        �Ͷ�m�$�H�p>�  ��������      ���������       �               ���       �� ?�  �       �������������������        �� ?�  �       @       ���      �         �����        �����  �XI$�H�m���I��       ���������       �         �      ���       �     ?         �������������������        �     ?         �       ��@               ������        �����  �|�  �������       �������        �         �      ���       ?��    �        A�����������?�������#�        ?��    �        A        ��       "          ����         ����m�$�H�~�  �������       ?�������        |         �      ���       ?��   �         �������������������G�         ?��   �         �        ����  ��D           ?����         |����  �[� H�l �I��       ?�������        >�         ��   ��p߀       ��   �        A�����������  ����  �� @       ��   �        A        �~  �    � @         ����         >�����  ���� ����p߀       �������        }�          ��   ����        ��   �        ������������  ���� � �       ��   �        �        �?  �    �         ����         }��m�$�H���� ������        �������        >�          �   ����        ��   �        ������������� ���� ?�!        ��   �        �        �� �    !           ����         >�����  �[`�H�m���I�        �������        @                 ��        ��� ��        ���������������������"        ��� ��        �        ����  ��@"           ��          @����  ��   �� ��        �������        �                  �         ��� ?��        ����������������������$         ��� ?��        �@        ����  ���$           ��          ����m�$�H��   ��  �         �������        �                  �         �����         �?���������������������(         �����         �         ����  �� (                        �����  �[l  H�l �I�         �����         �                   �         �����         ����������������������0         �����         �        ����  �� 0                        �����  ��   ��   �         �����         �                   �         �����         ����������������������          �����         �        � ���  ��                          ��m�$�H��   ��   �         �����          �                   �         �����         ���������������������          �����                 �                                    �����  �$�6�m�$�I#m��         �����          |                   �          �����         ?����������������������           �����         ?�        �                                    |����  �  ���   ���          �����          >                   �          ���          ����������������������           ���          �        �                                    >���m�$�H�  ���   ���          ���                              �          ���          ����������������������           ���          ��       �                                    ����  �$�6�m�$�I#m��          ���           �                  �           ?�           ���������������������            ?�           �@       �                                    �����  �  ���   ���           ?�            �                  �                        �?��������������������                         �        �                                    �I$�6�m�'  ���   ���                         �                  �                        ���������������������                         �       �                                    �   ���$�6�m�$�I#m��                         �                  �                         ���������������������                          �       �                                    �   ���  ���   ���                          �                  �                         ��������������������                                 �                                     �I$�6�m�'  ���   ���                          |                  �                         ?���������������������                          ?�       �                                     |   ���$�6�m�$�I#m��                          >                  �                         ���������������������                          �       �                                     >   ���  ���   ���                                            �                         ���������������������                          ��      �                                     I$�6�m�'  ���   ���                          �                 �                         ��������������������                          �@      �                                     �  ���$�6�m�$�I#m��                          �                 �                         �?�������������������                          �       �                                     �  ���  ���   ���                          �                 �                         ��������������������                          �      �                                     �$�6�m�'  ���   ���                          �                 �                          ��������������������                           �      �                                     �  ���$�6�m�$�I#m��                           �                 �                          �������������������                                 �                                      �  ���  ���   ���                           |                 �                          ?��������������������                           ?�      �                                      }$�6�m�'  ���   ���                           >                 �                          ��������������������                           �      �                                      >  ���$�6�m�$�I#m��                                            �                          ��������������������                           ��     �                                        ���  ���   ���                           �                �                          �������������������                           �@     �                                      ��6�m�'  ���   ���                           �                �                          �?������������������                           �      �                                      � ���$�6�m�$�I#m��                           �                �                          �������������������                           �     �                                      � ���  ���   ���                           �                �                           �������������������                            �     �                                      ��6�m�'  ���   ���                            �                �                           ������������������                                 �                                       � ���$�6�m�$�I#m��                            |                �                           ?�������������������                            ?�     �                                       | ���  ���   ���                            >                �                           �������������������                            �     �                                       >�6�m�'  ���   ���                                            �                           �������������������                            ��    �                                        ���$�6�m�$�I#m��                            �               �                           ������������������                            �@    �                                       ����  ���   ���                            �               �                           �?�����������������                            �     �                                       �6�m�'  ���   ���                            �               �                           ������������������                            �    �                                       ����[m�$�H�m�ܒI�                            �       �����  �                            ����������    ���                             �    �  �����                               ������������ �                             �         �   �                            ��������� � ���                                 �  ��?��                                �6�m�'�������� �                             |         0   �                            ?���������� 0 ���                             ?�    (�  �����                                |���[m�/�����ܒI�                             >    7         �                            ����������   ���                             �    H�  �����                                >���7�������� �                                 w     @   �                            ���������� @ ���                             ��   ��  �����                                I$�Hw�������� �                             �   �     @   �                            �������� @ ���                             �@  �  �����                                �   �[m�/�����ܒI�                             �  �     ��   �                            �?������� �� ���                             �   �  �|}��                                �  ��������� �                             �  �     ��   �                            �������� �� ���                             �  �  �x=��                                �$�K��������� �                             �  �     �B   �                             ����8���� �B ���                              �  8�  �x=��                                �  �[m�/����ܒI�                              �  �     ��   �                             ���x���� � ���                                x�  ��=��                                 �  ��������� �                              |       ��   �                             ?��������� � ���                              ?�   ��  ��}��                                 }$�_�������� �                              >  >     @   �                             ���������   ���                              �  A��  �����                                 >  >[m�/�����ܒI�                                }         �                             ��������� @ ���                              �� ���  �����                                   }�������� �                              � �         �                             �������   ���                              �@��  �����                                 ����������� �                              ��      0   �                             �?�	�����   ���                              � 	�  �����                                 ��[m�/�����ܒI�                              ��     �   �                             �������   ���                              �Ȁ  �����                                 ���������� �                              ��          �                              ��#�����    ���                               �#��  �����                                 ����������� �                               ��          �                              �G����    ���                               G�                                          ��[m�     ܒI�                               |p           �                              ?���������������                               ?� ��                                          |p��  ���� �                               >>�           �                              ��������������                               �A�                                          >����  ���� �                               }�           �                              ��������������                               ���                                          }�[m�$�H�m�ܒI�                               ��           �                              �������������                               �������������                                ��           �                               ���������������                              �                                            �                                             ���������������                               ��������������                              �@                                           �@                                            ��������������                               � �������������                               � �                                            � �                                            � �������������                                � �������������                               A                                             A                                              � �������������                                |                                              ?� �������������                               ?� �������������                                |                                               x                                              � �������������                               � �������������                                x                                               p                                              � �������������                               � �������������                                p                                               `                                              � �������������                               � �������������                                `                                               @                                              � �������������                               � �������������                                @                                                                                              � �������������                               � �������������                                                                                                                                � �������������                                � �������������                                                                                                                                  �������������                                  �������������                                                                                                                                  �������������                                  �������������                                                                                                                                  �������������                                  �������������                                                                                                                                  �������������                                  �������������                                                                                                                                  �������������                                  �������������                                                                                    ���������                                    ��        ��                                  ��        ��                                    ���������                                      ���������                                    ��        ��                                  ��        ��                                    ���������                                      ���������                                    ��        ��                                  ��        ��                                    ���������                                      ���������                                    ��        ��                                  ��        ��                                    ���������                                      ���������                                    ��        ��                                  ��        ��                                    ���������                                      ���������                                    ��        ��                                  ��        ��                                    ���������                                      ���������                                    ��        ��                                  ��        ��                                    ���������                                      ���������                                    ��        ��                                  ��        ��                                    ���������                                      ���������                                    ��        ��                                  ��        ��                                    ���������                                      ���������                                              @                                              @                                      ���������                                      ���������                                              @                                              @                                      ���������                                      ���������                                              @                                              @                                      ���������                                      ���������                                              @                                              @                                      ���������                                      ���������                                              @                                              @                                      ���������                                      ���������                                              @                                              @                                      ���������                                      ���������                                              @                                              @                                      ���������                                      ���������                                              @                                              @                                      ���������                                      ���������                                              @                                              @                                      ���������                                                                                      ���������                                      ���������                                                                                                                                      ���������                                      ���������                                                                                                                                      ���������                                      ���������                                                                                                                                      ���������                                      ���������                                                                                                                                      ���������                                      ���������                                                                                                                                      ���������                                      ���������                                                                                                                                      ���������                                      ���������                                                                                                                                      ���������                                      ���������                                                                                                                                      ���������                                      ���������                                                                                                                                      