�Sd  dN^r              x         l   �                           x         l   �                           x         l   �                           x         l   �                           � ��     �   �                           � ��     �   �                           � ��     �   �                           � ��     �   �                           � ��     �   �                           � ��     �   �                           � ��     �   �                           � ��     �   �                           ��<y����<���<�8                          ��<y����<���<�8                          ��<y����<���<�8                          ��<y����<���<�8                          y�f́���6f���3fٰ                          y�f́���6f���3fٰ                          y�f́���6f���3fٰ                          y�f́���6f���3fٰ                          �~�����6f�͘0fٰ                          �~�����6f�͘0fٰ                          �~�����6f�͘0fٰ                          �~�����6f�͘0fٰ                                                                                                                  �`�����6f�͘0fٰ                                                                                                                                                              ͛f́���6f�͘3fٰ                                                                                                                                                              x�<x�ٞ��<�͘<�3l                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            p                                 p        �                �                �                                                                                                �                �                �        �                �                �                                                                                             �                /�               �       �                /�               �       v                7`               v       r                '                r       �                /�               �       �                ?�               �       !                B               !                                                  q                G               q       �                o�               �        �               �                �                                                 > ��            ��>             > ��    ��            ��             ��    > C�            � >             > C�      �            �                 �    k F�            � k             k F�    *              ��*             *      w  'p            r w             w  'p    "                  "             "       �` 4             A�            �` 4    ]� }�            � �             ]� }�    �  8            0  c�            �  8    A                A             A      � "�            � *�            � "�    ~� #�            � >             ~� #�    �� �            � ɀ            �� �    H�  �            �               H�  �   �� 	�           �H  ��           �� 	�  �� π           ��  ��           �� π  �� ??�           �~ ��           �� ??�  �� �           �  ��           �� �  1i� T�`          � KF           1i� T�`  ?i� T��          �� K~           ?i� T��  0�� ?x`          ~ ��           0�� ?x`  0a� 0`           C           0a� 0`  n�@ ˰          �� <�           n�@ ˰  �@ ��          �� <�           �@ ��  N� �          �� �9           N� �  N@ Ð          �� <9           N@ Ð >�( ��[�        ��
8E��        >�( ��[��( ��y�        ��
8ǜ�        �( ��y�>�� ���        ��� �|��        >�� ����  #�I�        �� 8D��        �  #�I�k�  #�/�        �� 8B�`        k�  #�/�+�N  #�?�        �� 9�@        +�N  #�?�w?�� ���p        s�����w�        w?�� ���p#   #�'         2 � 8r@        #   #�' A� À,         �8�         A� À,]�N Ð=�        ��9ݠ        ]�N Ð=�c?�� ��0        3�� ��c`        c?�� ��0A  C�$         � 8A         A  C�$k�N C�n�        �� 9�`        k�N C�n��N  �?�        ��  9��        �N  �?�I?�� ��        ��� ��I         I?�� ��I   �$�        � �  8I         I   �$��@ �\           � 8�         �@ �\ ��0 #�}�        ��  8�܀        ��  �}�c� ?��0        1�� �|c`        c� ��0  �D           �  8@           �D K��  �<�        �� ���         K��P W�<��� �|�         ��  8��         �P S�|�w� �p        p�� 8w�        w  '�p   �          0 �  8 @            � 7�� �|         ���G�@        7�  %�| �� ~��         ��  �         �	  $�� ? �� w��        �� ߀~�        ? �� �� @ �         p �   @             � ��  G�        �� ��         �� �G�?�� ?��         ��p  p�         ?�� �� ~ �� 8��        �	 �?�        ~ � Fx�>               �                >       ��gP /w�        �����         ��w� Ow�}�U� �W�         ��P  Q�         }�U� MW� � �� ���        �
� ��?�        � �` 3��|             � @            |     ���H O_��        �����         ���TW��a�5� }w��        �P  P�         a�Etu��� �x {��        ����?�        � �� ���` �   �          @            `     �a��( V��0        ������         a�+� ���0a������0        �    �         a�:� ���0>�����        �.s�y�>�        >�0 g�  B "                                 1��� ��|`        �����         1����/�`1��� ���`        �(  ��         1���?|`>�< ���        �9�@	~`>�        >Dƃ�0
@ B `                        0   `9�S��+�`        �������@        9.K�`9������`        ��(  �/�@        9˚�:Μ`�v���        ��q�s�<�        <g �1��" B�@        ��                �@�I�-K��        �������         ���\_��+�~����        ��  @(L         k�^�~���{��y��        ��� �߼�        ��� /���H�  ���        ��  @         )�  ���)� \W7�        �������        �I� \�?���| ��]�        �P @R�        ��ru�}��� o���         ����9�         
�3��c��T �!(�         �@  @         �  � ��� ��          �߀���         ��� ��j ��x u��         �( @�         
��L��z� �?� ��          	�{��~@         G� o�  *A eP              @            A  @  [�� 8�h          ?�����          �� 9.x ��� ���           �  ��           �� �:� �w� ���          q� �s�          g� �0  *� BP              �            b � 0  Y�� y=h          ���݀         Y��y|�  m~� k��          
 �B          y|�i��  {�� ]�x          �<����          ��� �/�   � 
�             �@           	 � $�  ,�� zz�          ������          z�� �z�  �����|           J
 ��           ~�� �k�  ����_�          �����           1�� ]�`  �� 	��             ��           0�� `  ,�d ���          o���           ��z���  6�\ ��           � �           ��Z���  =�� ���          }�@��           G��8_  
�@ I@             �           �@ I   rt �u�          ���?o�          =ttqu�  }__���           %            ?\TQ��  w�����          �>���           �� �8�  
AH @                        @@ �  :rq�          ���~�           V�us�P  �^ׯ`           B� 
           ^�]׫�  s��y�          ?n ��           #t�9v   �@ &�                        $@ "   9:j�`          ���~�~           ::���  ������           � 
�           �*���  �{�{~`          ���>           q�|q�   � �)�                            !�   �9c�            =��>��           	�:��܀  ׯ�_            B             ׮��_�  ����            ��'/�            �qr�    R   H                          �  "X    ���            �����           �9�    ˯Ϯ�            ��
)            �)��    ���u�            	�p7�@           �y�    ("(�             �                 �    N��Ǩ            ��}��            �Eϸ   �ׇ^�             � (             ��G^�   �����            ��N_�            }8���    ) @�             �              i D�    WZ �h            }�-��           W���T    e�]X            Q@R            u���t    ~� ��            �/��            �{s�    Q              A               A     +�f�            �@g�            {�n�    ���j|             +x��             z�j�    �x ��            ��w             7z �`    0 b�             #               20 b`    )��<�            O��             ���:�    0��8�             ��             ���:�    ?����            ���             G���    ��8@             ��              ��:     O�            �D��            ?O�    O�             q�d�             ?O�    s����            �_��             ����     N@             0 D�              N�    R��            �e(�             WR�P    r�`             p�(�             _r��    ���            ?�"             #��       ��             0                 �     � �@            �b	�             � ��    ?�p��             x�	�             �p��    9��p             ��L             ��    � ��             @             � ��    �               �             )��    �!�             �b�             /�!�    ���              ��@             ���@    �               @             �     ��8              </��             ��:     ��?�            �o��             ��?     ���              /���             ���     ��              ,��             ��
     �9              \0c�             �9     �9�            �0c�             �=     ���              o���             ���     �	              L0`�             �	      � �              �               � �     � ��             ���              � �     ��              w��p             ��      h �              �	               h �     p f              w `             p f     p n              w �             p n     ���              {��p             ���     0 f              s `             0 f     �               �  �             �      �               �  �             �      ���              ���0             ���     �                �                �       ��             �@             ��     �             @@             �     ~��             �￰             ~��     @                               @       ��             �8�@             ��     ?���            ��L             ?���    �w�             ��             �w�     �                               �       ��            �@(             ��    �  �            �  *             �  �    9����            ����             9����    9   �            �               9   �   �p�@            P�T            �p�@   � ��            ��\            � ��    ��w�             ��             ��w�     �                P                �       ��@             <!?�             ��@    ��            8`              ��   y���             ����            y���                                             3�a@            0#8�            3�a@   � p!�            8            � p!�   ߏ�             ����            ߏ�                                              2`             0 &             2`    �@              X�            �@    ��r��            ?�+�            ��r��                                             D$!!�            4BB            D$!!�   V�             5`            V�   ����             ?�ʟ�            ����                                              "�p�             2/��            "�p�    #��             "=��            #��    � �              ��             � �      "                                 "       � �             0?��            � �    ��W�             8�}�            ��W�     ~ �              �
�              ~ �                                                 �؈�             =���            �؈�    ���             <�]�            ���     8�              �/�              8�                                                  ��!�             ~��             ��!�    ��Q�             ���            ��Q�     �               :�              �                                                  |��             ��;�             |��     ���             ��?�             ���      �                �               �                                                   ��              ��              ��     |�|             �pw�             |�|      ��               ��               ��                                                  ��              ��               ��      ���              ��              ���                      @                                                                  >��              �               >��      }��              ��               }��                                                                                          '�              �|               '�      ?��              ��               ?��                                                                                             ��               ��               ��      ��              ��               ��                                                                                              �                ?�               �       �                �               �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ? `  0~�          � �           0    ��                                                                                                                                     1�  0`           � �           1�    �                                                                                                                                      1�  0`           � �           00    �                                                                                                                                      1�o���`�         ��́�|p         0>s�����8                                                                                                                                    ?nٛ0|ݶ         �6o�v�         0;fm�`��l                                                                                                                                    0l��0`٘         ���f`         03fm����0                                                                                                                                    03lك0`ٌ         �6�f0         03fm� ��                                                                                                                                    03lٛ0`ٶ         �6m��f�         1�fm�`��l                                                                                                                                    0l���`ٜ         �����fp         3cͳ���8                                                                                                                                                                                                                            