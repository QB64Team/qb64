�}h  $# (                      0   8�            P   T@  8�     {��  ��  8�  8�     W�@  8�          ?��            L�@  sY�  L@  @�@  ��`  ��  L@  @�@  � `  ��� � 0  �   ��x ��� � x � x � | ��| � � � | ��� � � ��~ � | ��~ �� ��? � > ��? �  ?��     � �? >~�π   = p��=P�W�>�^��< �Bq��@B��(@=w�׀ �  ��  }����   |�� �, yw���    9�� X�D {���� �  � 	 {���� 	  ,��	 {���� 	  � 	 {���� 	  )� X�D {���� �  t�� �$ {w���    ��  }����    Bz	�@B�
(@=u�׀     =9���=Y�w�>���< '� �  >���   ��? � ? ��    ��~ �~ �� � > �q� �� �^~ �| �� �� ��� � � ��� ��� �� ��  ���  ��� ���  ���  ��  ��  ��  ��  �   _   ?��  _   �   �   �   �                                          