�l  �T�                                �    �     �                                                             �    �     �                                                             �    �     �                                                             �    �     �                                                             `  �     �                                                             `  �     �                                                             `  �     �                                                             `  �     �                                                                �     �                                                                �     �                                                                �     �                                                                �     �                                                             ��������<�8                                                            ��������<�8                                                            ��������<�8                                                            ��������<�8                                                            ��6l ��m�3fٰ                                                            ��6l ��m�3fٰ                                                            ��6l ��m�3fٰ                                                            ��6l ��m�3fٰ                                                             o�����m�0fٰ                                                             o�����m�0fٰ                                                             o�����m�0fٰ                                                             o�����m�0fٰ                                                                                                                                                                                                                   l���m�0fٰ                                                                                                                                                                                                                                                                                             l�6l���m�3fٰ                                                                                                                                                                                                                                                                                             Ǚ�����l�<�3l                                                                                                                                                                                                                                                                                                                                                                                                                                             0                                                0                                                                                                                                                                                                                                                      ,                                                ,                                                ,                        0                                                                                                                                                 `                        ^                        .                        ^                                                 .                        p                        N                                                .                                                                                                  ߀                       ^                        ߀                                                \                        a�                       �                        ;                        �                                                                         @�                       ��                       5                        ��                       @                        �                        À                       <�                       ~                        |                                                 0                       �                                               �                                               �                        �                       �                       9                        r                        �                                                 0                        �                       �                      z                       �                       �                       r                       ��                      y                        ��                      �                                                 `                       �                      ���                      ��                      ���                                             ��                      ��                      ��                      ��                     �                                                 �                       ��                     ��                     ���                     ��                     �                      ���                     ��                     ��                     ��|                     ��                                                ��                      ��                     ���                    ���                     ���                     �                     ���                     ���                    	��|                     ���                    ��                                              ��                     	���                    ����                    _���                    ����                      |                     ���                    9���                    ����                    � |<                    � |                                               |                     ��                    ���?�                   ����                    ���?�                     �                    ���                    ~���                   ���<                    1���                   ���                                              �                    ���                  7�����                  �����                  7�����                      <                    5���                   e���                  '�����                  ��<8                  /��<                                                <                    8���                   /���?                   |���                   /���?                      �                   ,x���                   0����                   <��8                   � |�                    |�                                               �                   `z |?�                   _� ���                  .~ ��                   _� ���                       8                   /z |?�                   q� |?��                  N^ ��                   � �8�                  .$ �8                                                8                    = ���                  �� ���                  ^� ���                  �� ���                                         \� ���                  a� ���                  �o ���                  ;R  <                  �R  <                                                                  @�  <?�                  ��  ?��                 5?  ?��                  ��  ?��                 @    �                  �=  <?�                  ý  <?��                 <�  ?�                  ~  ��                 |  ��                                           0    �                  �� ���                 7� ���                 �� ���                 7� ���                 �                      �� ���                 �>� ���                 9� ��                 r)   8p                 �	   8                                           0                       �  8��                 ?�  ?�|                 :�  ?��                 ?�  ?�|                      �                 r�  8��                 �  8��                 9�  ?�p                 ,	   �                 9	   �                                               �                 @  �                 �  ���                �  ��                 �  ���                      p                 @  �                 @  ��                �  ��                 �   �s�                �   �p                                                p                 @   ���                �   ���                 �   ���                �   ���                                       @   ���                @   ���                �   ��                 �   `                 �                                                                     �   �                 �   �x                 �   ��                 �   �x                      �                 �   �                 �   �                 �   �`                 
@   ��                 @   ��                                               �                 �   ��                 �   ��                 �   ��                 �   ��                       `                 �   ��                 �   ��                 �   ��                 
@    pg                 @    p`                                                `                 �    s�                 �    ��                �    �                 �    ��                                       �    s�                 �    s��                �    �                      �                                                                                      �    �                �    ��                �    ��                �    ��                                       �    �                �    �                �    ��                     �0                     �                                                                 �    ��                x    �<                �    ��                x    �<                 �      �                �    ��                �    ��                x    �0                �     `�                 �     `�                                          �      �                �     g�                x     �                �     �                x     �                 �      0                �     g�                �     g�                x     �                �     3                 �     0                                          �      0                 �     �                �     ��                �     �                �     ��                @                       �     �                �     ��                �     �                H     �                H                                               @                       �     ?�               �     ��                �     ��               �     ��                @                       �     ?�               �     ?�                �     ��               H      �0                H      �                                          @                       z      ��                �      �<                ~      ��                �      �<                        �                z      ��                �      ��                ^      �0                �      0�                $      0�                                                 �                z      3�                �      ?�                ~      ?�                �      ?�                        0                z      3�                �      3�                ^      ?�                �      3                $      0                                                 0                =      �                o      ��               ?      �                o      ��                                      =      �                }      ��               /      �                R      �                                                                                     =      ?�               o      ��               ?      ��               o      ��                                      =      ?�               }      ?�               /      ��               R       �0                      �                                                                �      ��               7�      �<               �      ��               7�      �<                       �               �      ��               >�      ��               �      �0               )       0�               	       0�                                                �               �      3�               7�      ?�               �      ?�               7�      ?�                       0               �      3�               >�      3�               �      ?�               )       3               	       0                                                0               @      �               �      ��              �      �               �      ��                                     @      �               @      ��              �      �               �      �              �                                                                     @      ?�              �      ��              �      ��              �      ��                                     @      ?�              @      ?�              �      ��              �       �0              �       �                                                               �       ��              �       �<              �       ��              �       �<                       �              �       ��              �       ��              �       �0              
@       0�              @       0�                                                �              �       3�              �       ?�              �       ?�              �       ?�                       0              �       3�              �       3�              �       ?�              
@       3              @       0                                                0              �       �              �       ��             �       �              �       ��                                    �       �              �       ��             �       �                      �                                                                                   �       ?�             �       ��             �       ��             �       ��                                    �       ?�             �       ?�             �       ��                      �0                      �                                                              �        ��             x        �<             �        ��             x        �<              �         �             �        ��             �        ��             x        �0             �        0�              �        0�                                       �         �             �        3�             x        ?�             �        ?�             x        ?�              �         0             �        3�             �        3�             x        ?�             �        3              �        0                                       �         0              �        �             �        ��             �        �             �        ��             @                       �        �             �        ��             �        �             H        �             H                                               @                       �        ?�            �        ��             �        ��            �        ��             @                       �        ?�            �        ?�             �        ��            H         �0             H         �                                       @                       z         ��             �         �<             ~         ��             �         �<                        �             z         ��             �         ��             ^         �0             �         0�             $         0�                                                 �             z         3�             �         ?�             ~         ?�             �         ?�                        0             z         3�             �         3�             ^         ?�             �         3             $         0                                                 0             =         �             o         ��            ?         �             o         ��                                   =         �             }         ��            /         �             R         �                                                                                  =         ?�            o         ��            ?         ��            o         ��                                   =         ?�            }         ?�            /         ��            R          �0                      �                                                             �         ��            7�         �<            �         ��            7�         �<                       �            �         ��            >�         ��            �         �0            )          0�            	          0�                                                �            �         3�          7�         ?�          �         ?�  �        7�         ?�                     0          �         3�  �        >�         3�   �        �         ?�   �        )          3   �        	          0                                                0   �        @         �?���        �         ��  �        �         �?���        �         ��  �                   ?���        @         �?���        @         �����        �         �  �        �         ����        �         ?���                        �                   ?���        @         ?� �        �         �����        �         �� �        �         ����                   @         @         ?�         @         ?����        �         �� �        �          ����        �          �@                                             @          �          π         �          ���        �          ��         �          ���                    �         �          π         �          �����        �          �  �        
@          0����        @          0�                                              �          �          9� X        �          ?���X        �          ?� X        �          ?���                    @         �          9�         �          9����        �          ?� �        
@          ���        @          @                                              @          �                    �          ���        �          �         �          ���                              �                    �          ���        �          � �                   ����                   �                                                           �          � �        �          ����        �          � �        �          ���                              �          �         �          ����        �          � �                    ���                                                                                �           /���        x           ���        �           /���        x           ���         �              �        �           /���        �           ��        x           /��        �           P          �                                                 �                      �           =         x           o         �           ?         x           o          �                    �           =         �           }  �        x           /  �        �           R  �         �                                              �                      �           =  �        �           o  �         �           ?  �        �           o  n         @             n         �           =  n        �           }  0         �           /  0        H           R  0         H                                                @                       �           =  s        �           o  s         �           ?  s        �           o           @                      �           =          �           }  �         �           /  �        H           R  �         H             `                        `         @             `         z           =  �         �           o  �         ~           ?  �         �           o �@                     �@        z           = �@        �           }   �        ^           /   �        �           R   �        $                                                                        z           =  �        �           o  �        ~           ?  �        �           o  <�                      <�        z           =  <�        �           }  �        ^           /  �        �           R  �        $             �                       �                      �        =           =  ;         o           o  ;         ?           ?  ;         o           o  �                     �        =           =  �        }           }           /           /           R           R                                                                               =           =  �        o           o  �        ?           ?  �        o           o  �                     �        =           =  �        }           }  8         /           /  8         R           R  8                                                                             �          =   �        7�          o   �        �          ?   �        7�          o  o�                     o�        �          =  o�        >�          }            �          /            )           R            	                                                                       �          =  0        7�          o  0        �          ?  0        7�          o  0                     0        �          =  0        >�          }  �        �          /  �        )           R  �        	                                                                    @          =  �        �          o  �        �          ?  �        �          o  �                     �        @          =  �        @          }           �          /           �          R           �                                                                   @          =  0        �          o  0        �          ?  0        �          o  �                     �        @          =  �        @          }           �          /           �          R           �                                                                   �          =  0        �          o  0        �          ?  0        �          o  �                     �        �          =  �        �          }           �          /           
@          R           @                                                                      �          =  �        �          o  �        �          ?  �        �          o  �                     �        �          =  �        �          }  8        �          /  8        
@          R  8        @                                                                �          =  �        �          o  �        �          ?  �        �          o  �                     �        �          =  �        �          }   �        �          /   �                   R   �                      �                        �                      �        �          =  �        �          o  �        �          ?  �        �          o  �                     �        �          =  �        �          }  �        �          /  �                   R  �                     �                       �                     �        �          =          x          o          �          ?          x          o  �         �            �        �          =  �        �          }           x          /           �          R            �                                                �                      �          =   s        x          o   s        �          ?   s        x          o   �         �             �        �          =   �        �          }   N        x          /   N        �          R   N         �             B                        B         �             B         �          =   �        �          o   �         �          ?   �        �          o   o         @             o         �          =   o        �          }   0         �          /   0        H          R   0         H                                                @                       �          =   `        �          o   `         �          ?   `        �          o   ~         @             ~         �          =   ~        �          }   �         �          /   �        H          R   �         H             `                        `         @             `         z          =            �          o            ~          ?            �          o                                 z          =           �          }   �         ^          /   �         �          R   �         $                                                                        z          =            �          o            ~          ?            �          o   ߀                      ߀        z          =   ߀        �          }            ^          /            �          R            $                                                                     =          =   �        o          o   �        ?          ?   �        o          o   /�                     /�        =          =   /�        }          }            /          /            R          R                                                                                =          =   �        o          o   �        ?          ?   �        o          o   �                     �        =          =   �        }          }            /          /            R          R                                                                                �         =   @        7�         o   @        �         ?   @        7�         o   �                     �        �         =   �        >�         }            �         /            )          R            	                                                                    �         =   @        7�         o   @        �         ?   @        7�         o   �                     �        �         =   �        >�         }            �         /            )          R            	                                                                    @         =   �        �         o   �        �         ?   �        �         o   �                     �        @         =   �        @         }            �         /            �         R            �                                                                   @         =   �        �         o   �        �         ?   �        �         o   �                     �        @         =   �        @         }            �         /            �         R            �                                                                   �         =   �        �         o   �        �         ?   �        �         o   �                     �        �         =   �        �         }   �        �         /   �        
@         R   �        @            �                       �                     �        �         =   �        �         o   �        �         ?   �        �         o   �                     �        �         =   �        �         }   �        �         /   �        
@         R   �        @             �                        �                      �        �         =   �        �         o   �        �         ?   �        �         o                                 �         =            �         }   �        �         /   �                  R   �                                                                            �         =   � �      �         o   �        �         ?   � �      �         o                          �      �         =    �      �         }   � �      �         /   �                  R   � �                     �                                             �      �         =   �      x         o   ��      �         ?   �      x         o   �       �                     �         =         �         }   ��      x         /   �      �         R   � �       �                                              �                     �         =    � 8      x         o   ��      �         ?    � 8      x         o   ��       �             �        �         =    �        �         }   ��      x         /    � 8      �         R   ��       �             �                        �         �             �         �         =     |      �         o    ���       �         ?     |      �         o    ��       @              8       �         =     8      �         }    ���       �         /    p |      H         R    ���       H              8                        8       @              8       �         =    �|      �         o   ��       �         ?    �|      �         o   ��       @             �(       �         =    �(      �         }   ���       �         /     |      H         R   ���       H             �(                        (       @             �(       z            � |       �           ���       ~            ��|       �           ���                     � 8       z            � 8       �           ���       ^             �|       �         ~  ����       $             ��8                        8                     � 8       z            � 8       �          ����       ~            ���8       �          ����                    �          z            �         �          �� �       ^             ��8       �          �����       $            ���                                              �          =          � �        o         �������       ?          ����       o         �������                 �           =          � �        }         ��� ��       /            ���       R         ������                  ���                                           �           =         >� � �       o        ����� �       ?         >���� �       o        ����� �                "�            =         "� � �       }        ��� � �       /          ��� �       R        �����                    ���                                             �            �          �          7�       �����          �        ?���          7�       �����                   ]              �        ]  �          >�       �� �          �        "���          )        ����           	          ?��                                                            �         �           7�       ����           �        ?��           7�       ����                    ]              �        ] �           >�       ���           �        *?��           )        ���            	         ?�                                                           `        �            �       ���            �       ?�            �       ���                     ]              `        ]�            `       ���            �       "?�            �       ��             �                                                                       �        >              �       ��             �       >              �       ��                      "              �        "              �       ��             �                     
@       ��             @                                                                       �                   ����������             �                   ����������             �                   �                   ����������             p                      ����������             �                                               �                      ���������               �       �              ����������              �       �               ��������               ���������               ���������              �     �              ���������               ���������                                        ��������                      �              ����������              ����������              ����������                                            �                     �              ����������              ���������>              ���������                                                                                      ����������               ����������               ����������                                                                                      ����������               ����������               ����������                                                                 ��������                ��������                ��������                ��������                                         ��������                ��������                ��������                                                                                                                                                                                                                                                                                                                                                                                                                �                       �                       �                                                                                                  �                       �                       �                                                                                                  ?�    `                  ?�    `                  ?�    `                  �����                  �����                  �����                  ;�                       ;�                       ;�                                                                                                  ?������                  ?������                  ?������                                                                                             ?������                  ?������                  ?������                                                                                             �    x                  �    x                  �    x                                                                                          �    h                  �    h                  �    h                                                                                                   <                        <                        <                                                                                                4                        4                        4                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ����                      |�0|�                    >c~>a�                                                                                                                                                                                                                                                  a��0                      f�0��                    cccca�                                                                                                                                                                                                                                                  c��0                      f�x��                    `cccs�                                                                                                                                                                                                                                                  c��0                      f�x��                    `cccs�                                                                                                                                                                                                                                                  �f�0                      |����                    `~c�                                                                                                                                                                                                                                                  f�0                      f����                    `ccc�                                                                                                                                                                                                                                                  ��0                      f����                    `cccm�                                                                                                                                                                                                                                                  6�0                      f����                    ccccm�                                                                                                                                                                                                                                                  6�0                      |��|�                    >cc>a�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         PP                   �
�   @     �         �
�    @       P                                                                                                                                                                                                                                        �P                   �    @     �         �     @       P                                                                                                                                                                                                                                        ��P                  �    @     �        �     @       P                                                                                                                                                                                                                                        ��P9c�<�8��c�          ��v9XN9 ��g��      ��v9XY��pq�3ӌ`                                                                                                                                                                                                                                      ��PE�YEE��Q          ��IdAE@	AH��       ��Ide"��� �TR�                                                                                                                                                                                                                                      �QPA�E�A�G�          
���I=DOA�	�OH���      
���I=DE"���'�W�@                                                                                                                                                                                                                                      �QPAQE A�$          
���IEDQA@	QH�@      
���IEDE"���(�T                                                                                                                                                                                                                                       �!PEQEE��Q          B��IEDQE 	QH��       B��IEDE"���(�TR�                                                                                                                                                                                                                                      �!P9�<�8��c�          B��I=DO9��G��      B��I=DE�qq�ӌ`                                                                                                                                                                                                                                      �                                   @                                                                                                                                                                                                                                                                  @     x                   �           �           �            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �                             �                      �                                                                                                                                                                                                                                                 �                      @      @               @      @                                                                                                                                                                                                                                                 �                      @      @               @      @                                                                                                                                                                                                                                             ,���,s��                `q��r�;@              `q��r�;@                                                                                                                                                                                                                                             ����(��J$                @�*(�(��@              @�*(�(��@                                                                                                                                                                                                                                             �"���"�K�                @�*(�/��@              @�*(�/��@                                                                                                                                                                                                                                             �"��H"�J                @�*(�($�@              @�*(�($�@                                                                                                                                                                                                                                             ����(��J$                @�*(�(��@              @�*(�(��@                                                                                                                                                                                                                                             "���"rI�                @q��r'$�@              @q��r'$�@                                                                                                                                                                                                                                                                                 @                        @                                                                                                                                                                                                                                                                                 �                        �                                                                                