��g  X  ��������������������������p��p��p��p��0��0��0��0������������������0��0��0��0� p� p� p� p� �� �� �� ������������������������������������������?��?��?��?��������������������������������������������������������������������� �     �    �    <    �    �    �                               �      @ �      �   `    1�    �    c�   A�    ǀ 8  �    �  p       �     < �     x � 0    �   `    1�    �    c�   A�    G� 8         0                                                   ��< '� �  >���   ��? � ? �� 