�gd  `�Oa                                                                                                                                                                                                                                                                                                                                                                                            "                                         "                                                                                  >                                         A                                         A                                         >                                                                                  ��                                        ��                                                                                 ��                                       @                                       @                                        ��                                       ��                                                                                                                       ��                                       ��                                       .                                       .                                       ��                                       ��                                       O                                       O                                       ��                                       px                                       ��                                       ��                                       px                                       �<                                       !�                                       !�                                       �<                                       =�                                       B?�                                       B#�                                       =�                                       {�                                       ���                                      �A��                                      {�                                       � �                                     ��@                                     ��@                                      �I�                                     � �                                     ��                                       |                                      ��                                     � �                                     #��                                     " >                                     ݀�                                     �  �                                     G��                                     D                                      �� �                                     p  x                                     ����                                     � �                                     w� x                                     �  <                                     !���                                     ! �                                     � <                                     =�                                       B?���                                     B  �                                     =��$                                     {�                                       �����                                    �@ ��                                    {��                                      �   �                                   ����@                                   �  �@                                    �� �                                   �   �                                   ����                                       |                                    �m�$��                                   �   �                                   #����                                   "   >                                   ��� �                                   �    �                                   G����                                   D                                      ���  �                                   p    x                                   ������                                   �   �                                   sm�$�x                                   �    <                                   !�����                                   !   �                                   ���  <                                   =�                                       B?�����                                   B    �                                   =���                                     {�                                       �������                                  �@   ��                                  {�m�$�                                   �     �                                 ������@                                 �    �@                                  ���  �                                 �     �                                 ������                                       |                                  ����  �                                 �     �                                 #������                                 "     >                                 ��m�$�A�                                 �      �                                 G������                                 D                                      ����   �                                 p      x                                 ��������                                 �     �                                 w���   x                                 �      <                                 !�������                                 !     �                                 ��m�$�H<                                 =�                                       B?�������                                 B      �                                 =����                                    {�                                       ���������                                �@     ��                                {����                                    �       �                               ��������@                               �      �@                                �6�m�$�H�                               �       �                               ��������                                       |                                �����  ��                               �       �                               #��������                               "       >                               �����  ��                               �        �                               G��������                               D                                      ���m�$�H��                               p        x                               ����������                               �       �                               w����  �x                               �        <                               !���������                               !       �                               �����  �<                               =�                          p            B?���������                               B        �                  p            =�I$�6�m�$                               {�                          �            �����������                              �@       ��                 �            {�   ���                                �         �                �           ����������@                           �        �@                �            �`   ��� �                           �         �                �           ����������                Q                    |                 �           �rI$�6�m�$��               q           �         �               �           #����������              #           "         >               �           ��   ��� �              #           �          �             ?� �           G����������                         D                      ?� �           ��   ���  �                         p          x             �  �           ������������                         �         �             �  �           srI$�6�m�$�x                         �          <             �� p           !�����������              �           !         �             �� p           ��   ���  <              �           =�                       ��8             B?�����������                        B          �             ��8             =��   ���               
           {�  �                    ��  �         ������������                     �@  �      ��            ��  �         {�rI��6�m�$�                      �  d       �           ������        ������������@             4         � �       �@           ������         ��� ���  �            ���4         �  �       �            �����        �����������              �@          �       |             �����        ���� ���  �             ����@        �  �       �            ���?�        #������������            �/�         "         >            ���?�        ��rO��6�m�$�A�            �?���         �  �       �            ?� 8 ?�        G����������           ��:Ā        D  ��                  ?�   >�        ��������   �           ��ŀ        p  ��       x               ?�        �������������           ��?�@        �  �      �                >x        w�������   x           ��?��        �  ��       <             �  ?�        !������������           �"?��       !  �      �             �  >x        ��rO��6�m�$�H<           �"?���       =�  �                   � ��        B?������������           �&�@@       B   �      �            �  ?�        =�������              �&D@@       {�  �                    � ��        ��������������          �L�?�         �@  �      ��            �  �        {�������              ��8          �           �            � ��       ��������������@         ���T�        �          �@            �  ��        �6�rO'�6�m�$�I�         ���Tx�        �   �        �             � ��       ��������������          ��oH��                   |              � ��       ����� ���   �         ��oL��0       �    �        �          p   �8       #�������������          ��Ο��       "   �        >          p     �8       ����� ���   �          �x�Μ��       �    p         �          � �   x       G�������������          �?���       D    �                  �      x       ���rI��6�m�$�I �          �0|��       p              x          � �          ����������������          �?��g        �             �          �            w���   ���    x          '�"<�g       �              <         �p�  �       !���������������          �����        !             �         �    �       ����   ���    <         ��?��       =�                       ���  �       B?���������������          ����?�        B              �         �    �       =Ͷ�rI$�6�m�$�I          ��>�?�       {�                       ���  �       �����������������         �������      �@             ��        �     �       {����   ���            �'�����      �               �          �   �      ����������������@        ���� �     �              �@               �       ����   ���   �        �C����     �               �         p    ��     ����������������          ����2�                     |               ��     �m��rI$�6�m�$�I#�        ����2��     �               �             ��     #����������������         �����8>      "               >              ��     �����   ���   ��        �����8>�     �                �            > ��     G����������������         �����<      D                             ��     �����   ���   ��        �����<�     p                x           >   p     ������������������        �����ÿ��     �               �              p     t�I$���m�$�H�m�ܐx        �����˿��     �                <           >>  p     !�����������������        ����?���      !               �           >   p     �   ����  ���� <        �������p     =�                        8 �  8     B?�����������������         �澈       B                �        8 @   8     =�   ����  ����         8�f>� 8     �                        8 �  �8     a������������������        �����       a@               ��       8      8     ��I$���m�$�H�m�ܒ        8d��� 8                      �       8 � � 8     p������������������@        ������      p�                �@       8     8     x   ����  ���� �       8�����8     �                �       x�> � <     x�����������������         �������      x@                |        x �>  @ <     �   ����  ���� �       x�����G�<     �                �         � �      |?�����������������       ���~����      |                 >         @  �      ܒI$���m�$�H�m�ܒA�       ��������     �                 �       p �  �      ~�����������������      ����������     ~                       p �   @      �   ����  ����  �      �������G��      �                 x       p �  �      ������������������       ��g�����                     �       p              �   ����  ����  x      p�g����      x                 <       p �  �      �������������������       {d�G���      �                �       p @           x�I$���m�$�H�m�ܒH<      p{�>G��       <                        �           �������������������       �C��D��=�     �                �       p            <   ����  ����         �C��D��=�                              �   ��      ��������������������      ���<@7�     �                ��      p   ��          ����  ����         ���4@7�                       �      �   �      �������������������@      ���΀'�     ��                �@      p   �       I$���m�$�H�m�ܒI�      ���΀'�      �                �      � �  ��      ������������������       �7��� �     �@                |       p    ��       �  ����  ����  �      �7��@�      �                �     � � ��      �?�����������������     �w���~  C     �                 >      p    ��       �  ����  ����  �     �w��~  _      �                 �     � � �� ?     ������������������     ���_�~       �                      x    �� <      �I$���m�$�H�m�ܒI �     ������ ?       �                 x     � �8�� ;     �������������������     �'���� ��     �                �      8  @ �� <       �  ����  ����   x     �'�G��.��?       x                 <     ���|�� ;     ��������������������     �?_��  `     ��                �      8�  �� <       x  ����  ����   <     �<��� `?       <                      ���|�� ;     ��������������������     �����     ��                �      8� �� <       <I$���m�$�H�m�ܒI$     ����?                             ���|�� s     ���������������������    ���n�      ��                ��     � ( �� |         ����  ����        ��:�                         �    �� 8� s     ��������������������@    �0�> 8     ���                �@     �  � |         ����  ����   �    �0� 8       �                �    ��   ?� �     �������������������     �"��@<     ��@                |      �   ?� �       �$���m�$�H�m�ܒI$��    �"��@<�       �                �    �       �     ��?�����������������    ���`�     ��                 >            �       � ����  ����   �    ���`��       �                 �    �       �     �������������������    �����      ��                            �       � ����  ����    �    ������        �                 x    �       �     ?��������������������    �����      ?��                �            �        �$���m�$�H�m�ܒI$�x    ������        x                 <    ��     �     ���������������������    ���?�      ���                �     �      �        x ����  ����   <    ����7��        <                     ��           ���������������������    �~?�      ���                �     �      �        < ����  ����       ��~?��                              �� �        ����������������������    ���      ���                ��    � �   �        $���m�$�H�m�ܒI$�     �����                         �    �� �        ���������������������@    �  ��      ����                �@     � �   �         ����  ����   �    �� ���        �                �    �� �   x     ��������������������     �� ��      ���@                |      < �   �        �����  ����   ��    �� ���        �                �    �� �   �      ���?�����������������    �� ���        ���                 >     > �   ��        �rI$�6�m�$�I#m��rA�    �� ��� ��        �                 �    � �  �      �������������������    �          ��                      �  ��        ��   ���   ���� �    �  ��         �                 x    ���  �      ?��������������������    �  
        ?��                �     ��  ��         ��   ���   ���� x    �� 
��         x                 <    ���  �      ���������������������    �  �        ���                �     ��  ��         {rI$�6�m�$�I#m��rH<    �� ���         <                     ?��    > 8      ���������������������    ?�  	  8      ���                �     �    ?��         =�   ���   ����     ?�� 	?��                              ?�|    | x      ����������������������   ?�     x      ���                ��    �    ��         �   ���   ����     ?��  ��                          �   ?�?   � x      ���������������������@   ?�      x      ����                �@    �   ���         rI$�6�m�$�I#m��rI�   ?��  ���         �                �   ��  ?� �      ��������������������    �       �      ���@                |     ��  ?��          �   ���   ���� �   ���  ?���         �                �   ���  ?���       ���?�����������������   ��    ��       ���                 >     �  ?�          �   ���   ���� �   ���  ?���         �                 �   ������       �������������������   ��    �       ��                     �����          �I$�6�m�$�I#m��rI �   ��������          �                 x   �|?���|�       ?��������������������   �|    |�       ?��                �     �������           �   ���   ����  x   ���������          x                 <   �������       ���������������������   ��   ��       ���                �     p�����           x   ���   ����  <   ���������          <                    ���  ?��       ���������������������   ���  ?��       ���                �     <����           <I$�6�m�$�I#m��rI$   ���������                              ����� �       ����������������������  ����� �       ���                ��     ���              ���   ����     ���������                           �  ����� �       ���������������������@  ����� �       ����                �@    �  ?��              ���   ����  �  ���������          �                �  �� �  ?        ��������������������   �� �  ?        ���@                |     �����           �$�6�m�$�I#m��rI$��  ��������           �                �   ��     ~         ���?�����������������   ��     ~         ���                 >    ������           �  ���   ����  �   ��������           �                 �   �    �         �������������������   �    �         ��                     �����            �  ���   ����   �   �������            �                 x   ��   �         ?��������������������   ��   �         ?��                �     ����             �$�6�m�$�I#m��rI$�x   �������            x                 <   ?��   �         ���������������������   ?��   �         ���                �     ����             x  ���   ����   <   ?�������            <                    ��   �         ���������������������   ��   �         ���                �     ����             <  ���   ����      �������                                ��   ��         ����������������������  ��   ��         ���                ��    ���              $�6�m�$�I#m��rI$�   �������                             �  ��� ��         ���������������������@  ��� ��         ����                �@     ?��                ���   ����   �  �������            �                �  ��� �          ��������������������   ��� �          ���@                |      ��              � ���   ����   �  ������             �                �   ������           ���?�����������������   ������           ���                 >                      Ē6�m�$�I#m��rI$��   ������             �                 �   ?�����           �������������������   ?�����           ��                                      � ���   ����   `�   ?�����              �                 x   �����           ?��������������������   �����           ?��                �                       � ���   ����   px   �����              x                 <   �����           ���������������������   �����           ���                �                       x�6�m�$�I#m��rI$�0<   �����              <                    ����            ���������������������   ����            ���                �                       < ���   ����   |   ����                                    ?���            ����������������������   ?���            ���                ��                       ���   ����   ~    ?���                                �   ���            ���������������������@   ���            ����                �@                      m�$�H�m�ܒI$���m��   ���               �                �    �             ��������������������     �             ���@                |                       ��  ����   �����    �                �                �                    ���?�����������������                    ���                 >                      ߀  ����   �����                      �                 �                    �������������������                    ��                                      ��$�H�m�ܒI$���m� �                       �                 x                    ?��������������������                    ?��                �                       ��  ����   ���� x                       x                 <                    ���������������������                    ���                �                       {�  ����   ���� <                       <                                     ���������������������                    ���                �                       =�$�H�m�ܒI$���m�$                                                            ����������������������                   ���                ��                      �  ����   ����                                         �                   ���������������������@                   ����                �@                         ����   ���� �                      �                �                   ��������������������                    ���@                |                       �$�H�m�ܒI$���m�$��                      �                �                    ���?�����������������                    ���                 >                      �  ����   ���� �                      �                 �                    �������������������                    ��                                      �  ����   ����  �                       �                 x                    ?��������������������                    ?��                �                       �$�H�m�ܒI$���m�$�x                       x                 <                    ���������������������                    ���                �                       x  ����   ����  <                       <                                     ���������������������                    ���                �                       <  ����   ����                                                              ����������������������                   ���                ��                      $�H�m�ܒI$���m�$�                                        �                   ���������������������@                   ����                �@                        ����   ����  �                      �                �                   ��������������������                    ���@                |                       � ����   ����  �                      �                �                    ���?�����������������                    ���                 >                      ĒH�m�ܒI$���m�$�A�                      �                 �                    �������������������                    ��                                      � ����   ����   �                       �                 x                    ?��������������������                    ?��                �                       � ����   ����   x                       x                 <                    ���������������������                    ���                �                       x�H�m�ܒI$���m�$�H<                       <                                     ���������������������                    ���                �                       < ����   ����                                                               ����������������������                   ���                ��                       ����   ����                                           �                   ���������������������@                   ����                �@                      H�m�ܒI$���m�$�H�                      �                �                   ��������������������                    ���@                |                       �����   ����  ��                      �                �                    ���?�����������������                    ���                 >                      �����   ����  ��                      �                 �                    �������������������                    ��                                      �H�m�ܒI$���m�$�H��                       �                 x                    ?��������������������                    ?��                �                       �����   ����  �x                       x                 <                    ���������������������                    ���                �                       x����   ����  �<                       <                                     ���������������������                    ���                �                       =�$�I#m��rI$�6�m�$                                                            ����������������������                   ���                ��                      �   ����   ���                                         �                   ���������������������@                   ����                �@                      ~   ����   ��� �                      �                �                   ��������������������                    ���@                |                       �$�I#m��rI$�6�m�$��                      �                �                    ���?�����������������                    ���                 >                      �   ����   ��� �                      �                 �                    �������������������                    ��                                      �   ����   ���  �                       �                 x                    ?��������������������                    ?��                �                       �$�I#m��rI$�6�m�$�x                       x                 <                    ���������������������                    ���                �                       z   ����   ���  <                       <                                     ���������������������                    ���                �                       <   ����   ���                                                              ����������������������                   ���                ��                      $�I#m��rI$�6�m�$�                                        �                   ���������������������@                   ����                �@                         ����   ���  �                      �                �                   ��������������������                    ���@                |                       �  ����   ���  �                      �                �                    ���?�����������������                    ���                 >                      ĒI#m��rI$�6�m�$�A�                      �                 �                    �������������������                    ��                                      �  ����   ���   �                       �                 x                    ?��������������������                    ?��                �                       �  ����   ���   x                       x                 <                    ���������������������                    ���                �                       x�I#m��rI$�6�m�$�H<                       <                                     ���������������������                    ���                �                       <  ����   ���                                                               ����������������������                   ���                ��                        ����   ���                                           �                   ���������������������@                   ����                �@                      I#m��rI$�6�m�$�I�                      �                �                   ��������������������                    ���@                |                       � ����   ���   �                      �                �                    ���?�����������������                    ���                 >                      � ����   ���   �                      �                 �                    �������������������                    ��                                      �I#m��rI$�6�m�$�I �                       �                 x                    ?��������������������                    ?��                �                       � ����   ���    x                       x                 <                    ���������������������                    ���                �                       x ����   ���    <                       <                                     ���������������������                    ���                �                       <I#m��rI$�6�m�$�I                                                             ����������������������                   ���                ��                       ����   ���                                           �                   ���������������������@                   ����                �@                       ����   ���   �                      �                �                   ��������������������                    ���@                |                       �#m��rI$�6�m�$�I#�                      �                �                    ���?�����������������                    ���                 >                      �����   ���   ��                      �                 �                    �������������������                    ��                                      �����   ���   ��                       �                 x                    ?��������������������                    ?��                �                       �ܒI$���m�$�H�m�ܐx                       x                 <                    ���������������������                    ���                �                       {�   ����  ���� <                       <                                     ���������������������                    ���                �                       =�   ����  ����                                                             ����������������������                   ���                ��                      ܒI$���m�$�H�m�ܒ                                        �                   ���������������������@                   ����                �@                      x   ����  ���� �                      �                �                   ��������������������                    ���@                |                       �   ����  ���� �                      �                �                    ���?�����������������                    ���                 >                      ܒI$���m�$�H�m�ܒA�                      �                 �                    �������������������                    ��                                      �   ����  ����  �                       �                 x                    ?��������������������                    ?��                �                       �   ����  ����  x                       x                 <                    ���������������������                    ���                �                       x�I$���m�$�H�m�ܒH<                       <                                     ���������������������                    ���                �                       <   ����  ����                                                              ����������������������                   ���                ��                         ����  ����                                          �                   ���������������������@                   ����                �@                      I$���m�$�H�m�ܒI�                      �                �                   ��������������������                    ���@                |                       �  ����  ����  �                      �                �                    ���?�����������������                    ���                 >                      �  ����  ����  �                      �                 �                    �������������������                    ��                                      �I$���m�$�H�m�ܒI �                       �                 x                    ?��������������������                    ?��                �                       �  ����  ����   x                       x                 <                    ���������������������                    ���                �                       x  ����  ����   <                       <                                     ���������������������                    ���                �                       <I$���m�$�H�m�ܒI$                                                            ����������������������                   ���                ��                        ����  ����                   �                      �                   ���������������������@               �  ����                �@                        ����  ����   �               �     �                �                   ��������������������                �  ���@                |                       �$���m�$�H�m�ܒI$��               �     �                �              �   ���?�����������������               �   ���                 >              �     � ����  ����   �               �     �                 �             D   �������������������               p   ��                             �     � ����  ����    �            |  �      �                 x               �   ?��������������������            |  �   ?��                �               �      �$���m�$�H�m�ܒI$�x            �  �      x                 <             0    ���������������������            �  �   ���                �             0       x ����  ����   <           �  �      <                              0    ���������������������           �  �   ���                �             0       < ����  ����              ��@�                                    8b   ����������������������          ��@�   ���                ��            8b      $���m�$�H�m�ܒI$�           ���                         �            8D   ���������������������@          ���     ����                �@           (8D       ����  ����   �          ��@       �                �          @<H   ��������������������           ǀ@    ���@                |           x<H      �����  ����   ��          ��ǯ ?�    �                �            <8P�   ���?�����������������          ǃǯ ?�  ���                 >           8?���     �rI$�6�m�$�I#m��rA�          ��Ϯ �    �                 �            <0Q��   �������������������          ��Ϯ �  ��                            ����     ��   ���   ���� �          �C V ��     �                 x           �0i�   ?��������������������          �C  ��  ?��                �           �0?�      ��   ���   ���� x           �� � ��     x                 <           ~0��   ���������������������           ��   ��  ���                �          �0	�      {rI$�6�m�$�I#m��rH<           |  @ ��     <                           �~pH�	   ���������������������           |    ��  ���                �          �~p�      =�   ���   ����             �  ��                                O�|p��   ����������������������           �  ��  ���                ��         O�|p��     �   ���   ����             � ��                      �         o�8<�  ���������������������@           �  ��  ����                �@         o�8<�q     rI$�6�m�$�I#m��rI�           � �     �                �         /�93���   ��������������������            �  �  ���@                |          /�83���      �   ���   ���� �           � ?�     �                �        ��81Q�     ���?�����������������           � ?�   ���                 >        ��81Q�       �   ���   ���� �           � �     �                 �        ���q#     �������������������           � �   ��                        ���q3g �     �I$�6�m�$�I#m��rI �        �    �      �                 x         ?���:~7    ?��������������������        �     �   ?��                �         ?���:r7�      �   ���   ����  x        � >   �      x                 <         ���<pn    ���������������������        �     �   ���                �         ���<po�      x   ���   ����  <        �     x      <                          ���4a�    ���������������������        `     x   ���                �         ����4a�x      <I$�6�m�$�I#m��rI$        ��   <                                �����    ����������������������       �    <   ���                ��       >����<         ���   ����          ��                          �        �����`    ���������������������@       �       ����                �@       ����`         ���   ����  �       �>   ?�      �                �        ���#�J~   ��������������������         �    ?�   ���@                |        ���#�J~      �$�6�m�$�I#m��rI$��        �   ?�      �                �       ����/�@    ���?�����������������              ;�    ���                 >       ���/�D      �  ���   ����  �       �    ?�      �                 �        ǿ�?��`    �������������������             ?�    ��                       ~��?��g      �  ���   ����   �       8    p �      �                 x        ������    ?��������������������       8      �   ?��                �       8�������      �$�6�m�$�I#m��rI$�x       8    � �      x                 <        ?�������    ���������������������       8      �   ���                �       8?�������      x  ���   ����   <       p   p�  �      <                        ������    ���������������������       p   p   �   ���                �       w����'.���      <  ���   ����          p   ��  !�                              ��� ���    ����������������������      p   �   !�   ���                ��      w��� ���      $�6�m�$�I#m��rI$�       � �p  p�                       �      ��� |�     ���������������������@      � �   p�   ����                �@      ���� � �        ���   ����   �      � �� � �      �                �       ��S���     ��������������������       �  �    �   ���@                |       �}�:S��x �      � ���   ����   �      � �� � �      �                �       ��#����     ���?�����������������      � A�    �    ���                 >      ��:#��?��      Ē6�m�$�I#m��rI$��     �@�� � �      �                 �       �����     �������������������     �@ �   �    ��                     �;����      � ���   ����   `�        �p � p       �                 x     �������     ?��������������������         p � p    ?��                �     �;�����p       � ���   ����   px     � �  � p       x                 <     ������     ���������������������     � @    p    ���                �     ��;���p       x�6�m�$�I#m��rI$�0<     � �  � 0       <                      ���������    ���������������������     �        0    ���                �     ���y���?��       < ���   ����   |     �    � 0                             ����� @    ����������������������    �       0    ���                ��    	�����| p        ���   ����   ~     �    t|  8                        �    ����� H    ���������������������@    �    |  0    ����                �@    ������ x       m�$�H�m�ܒI$���m��    �    .�  x       �                �     ��� ��    ��������������������     �    �  p    ���@                |     ���� ��x       ��  ����   �����    �p   �  x       �               �     ��: �     ���?�����������������    �p   �  p     ���                >    ���: �x       ߀  ����   �����    � � �� x       �            �    �     ����      �������������������    �    �� p     ��           �       ���x�!x       ��$�H�m�ܒI$���m� �    � � �� |        �            @    x    �����D      ?�������������������    �    �� p     ?��           �   �    ���?��D |        ��  ����   ���� x    � � �� �        x                 <    ���� <      ���������������?�����    �    �� �     ���           �   �    �����8< �        {�  ����   ���� <    � ���� �        <                x     ������      ��������������������     �   �� �     ���           �   �    ����� �        =�$�H�m�ܒI$���m�$x    ����� �                        �     8��� �     �������������������     �   �� �     ���           ?�       �8��8��        �  ����   ?���� �    ������ �                       �     p��XD?�     �������������������     �� @�� �     ����          �       �p>NHD?��           ����   �����    ����;���        �              �    �r?��|@�     ������������������2     p� ����     ���@          ��   2    �r<x�D@��        �$�H�m�ܒI$���m�#�    �� �� �        �              �    ����X �@      ���?���������� ����b     p� @� �      ���          ��   b    ���XH �A�        �  ����  ������    �    � �        �            �  <    ���A �@      ������������  �����     8    � �      ��         ���  �    ���A �C�        �  ����  �����<    �     | �         �            @  |    �w�A��       ?������������  ���     8     | �      ?��         ���  !�    ��A��#�         �$�H�m�ܒI'���m�|    �                x               <�    � w��G��       �������������  ?���            �      ���         ���  C    � w��G���         x  ����  �����<�    �                <              y�    � G��G�        �������������  ���            �      ���         ���  �    � G��G� �         <  ����  �����y�    �                              ��    � ��@��       �������������  ��            �      ���         ?���     � ��@���         $�H�m�ܒI?���m���    �                         �   ��    � 9�P��       ������������π ?��            �      ����        p��     � 9�P���           ����  �������    ��     <         �        0` @ ��    � 8S��       ������������` ��0     �     ?�      ���@        ϟ�� 0    ��8S��?�         � ����  ��������    �� �   x8         �        @ � ��    �  0G�8 8       ���?��������@ ���`     � �   �       ���        ���  `    �� 0W�8�         ĒH�m�ܒI����mǟ�    �� �  �8         �        �  ?�    �   o� 8       ���������� ����      � �  ��       ��       ���  �    ��  o�	��         � ���� ������?�    �� �  �8          �        �  �    �  "n  8       ?���������� ���      � �  ��       ?��       ���  !�    �� "n��          � ���� �������    �� �  �p          x         <��    ��   ,  p       ��������������       | �  ��       ���       ���  C     ��   ,��          x�H�m�ܒO����m���    �� �  �p          <        �  y��    ��   (  p       ���������������       > �  ��       ���       �{�  �     ��   (��          < ���� �����y��    �π   > p                  �  ���    �� 0 "  p       ��������������       ?�   ?��       ���       ?�{�      ���0 "?��           ���� ?��������     ���    � �                  �  ���     ��   $  �       ������������?��       �    ��        ����      �{�       ���  $���          H�m�ܒ����m���     ���   ��          �       @ ���     ��   8 �       ������������0       �   ��        ���@      ���� 0      ���  8���          ����� ���������     ���   ��          �        � ���     ��   0  �        ���?������ ����`       �   ��         ���      ���  `      ���  0���          ��������������     ��  � �          �        	  ?��     �      �        �������� �	����       ��  ���         ��     ���  �      ���  ����          �H�m�ܓ�����o?��     ��  ��           �          ��     �     �        ?�������� @���       ��  ���         ?��     ���  !�      ���  ����           �������������     ��� �x�           x        d  <���     ��    x�        ��������� 0���         ?� ���         ���     ���  C       ��� ����           x�������������     ?��������           <       �  y���     ?��   ��        ��������� ���         �����         ���     ���  �        ?���������           =�$�I#���I$y���     ?�<����                     ��߀     ?�<   ��        ���������  ��  @      ������         ���     ?���   @     ?���������           �   ����  ��߀     ��  �                       ���      ��  �          ���������  ?�� P�       �����         ����    ���  P�     ��������            ~   ���� ���      ��� � >            �       @ ��v      ��� � >         �������   ��0 �        |����         ���@    ��� 0 �      ��������            �$�I#���I#��v      ����  ~            �       � ���      ����  ~          ���?�����  ���`        ?�  ���          ���     ?��  `      ��������            �   ���� ���      ����  �            �        ?��      ����  �          ������� ����        � ��           ��    ��  �      ��������            �   ���� ?��      ��    �             �        ��      ��    �          ?������� ���        �����           ?��    ��  !�      ��������             �$�I#o��rI��      ��    �             x        <���      ��    �          �������� ���  �       �����           ���    ��  C  �     ��������             z   ���� <���      ��    �             <        y����     ��    �          �������� ���  @       �����           ���    ��  �  @     ��������             <   ���� y����      ���   ?�                     �����      ���   ?�          �������� ��            ����           ���    ��           ��������             $�I#m��rH�����      ��   �                     �����      ��   �          �������� ?�� @         ?����           ����    ��  @       �������                ���������      ?��  ��             �     @ ����      ?��  ��          ������� ��0 �         ���            ���@    � 0 �       ?�������             �  �������      ��  �              �     � �����      ��  �            ���?��������`           ���             ���     ?  `        ������              ĒI#m��rG�����      �����              �      ?����      �����            �����������           �              ��      �        ������              �  ����?����      ������               �      ����      ������            ?����������                           ?��      !�        ������               �  ��������       ������               x      <�����       ������            �����������   
                         ���       C   
       ������               x�I#m��r<�����       �����               <       y�����       �����            �����������                            ���       �          �����               <  ����y�����       ����                       ������       ����             ����������    "                         ���          "       ����                  ����������       ����                      ������       ����             ���������� @  B                         ����      @  B       ����                I#m��q������        ����                �     ����|        ����             ���������0 �  �                         ���@     0 �  �        ����                � ��������|        ��                 �     ������        ��               ���?������`                            ���      `          ��                 � ���������        ��                 �     ?�����        ��               ���������                            ��     �          ��                 �I#m��o?�����                             �     �����                          ?��������                            ?��     !�                               � ���������                             x     <������                          ���������                             ���     C                                x ����������                             <     y������                          ���������                             ���     �                                <I#m��y������                                  �������                          ��������                                ���                                        ����������                                 �������                          �������� @  @@                          ����    @  @@                              ����������                             �   ����                           �������0 �  ��                          ���@   0 �  ��                             �#m������                              �   ������                            ���?����`                              ���    `                                ����������                              �   ?�����                            �������                              ��   �                                ����?�����                               �   �����                            ?������                              ?��   !�                                 �ܒI�����                               x   <������                            �������                               ���   C                                  {�  <������                               <   y������                            �������                               ���   �                                  =�  y������                                  �������                            ������                                  ���                                       ܒH�������                                 �������                            ������ @  @@                            ����  @  @@                               x �������                               � ����                             �����0 �  ��                            ���@ 0 �  ��                               � ����                                � ������                              ���?��`                                ���  `                                  ܒG������                                � ?�����                              �����                                �� �                                  � ?�����                                 � �����                              ?����                                ?�� !�                                   � �����                                 x <������                              �����                                 ��� C                                    x�<������                                 < y������                              �����                                 ��� �                                    < y������                                  �������                              ����                                    ���                                        �������                                 �������                              ���� @  @@                              ���� @  @@                                 �������                                 �����                               ���|0 �  ��                              ���D0 �  ��                                 �����                                  ǟ�����                                ���8`                                  ���(`                                    ǟ�����                                  �?�����                                ���                                  ���                                    �?�����                                   ������                                ?���                                  ?���                                     ������                                   |������                                ���                                   ���                                      |������                                   9������                                ���                                   ���                                      9������                                   ������                                ���                                     ���                                        ������                                   ������                                ���   @@                                ���   @@                                   ������                                   ���                                 ��� � ��                                ��� � ��                                   ���                                    ��?��                                  ��� �                                  ��� �                                    ��?��                                    ����                                  �� �                                  �� �                                    ����                                    ����                                  ?�� �                                  ?�� �                                    ����                                    ����                                  �� �                                  �� �                                    ����                                    ����                                  �� '�                                  �� '�                                    ����                                    ����                                  �� C�                                    �� C�                                      ����                                    �  ��                                  �� ��@@                                  �� ��@@                                    �  ��                                    �                                     �� ���                                  �� ���                                    �                                       �  ~                                    �� �                                    �� �                                     �  ~                                     �  |                                    � ?�                                    � ?�                                     �  |                                     �  x                                    ?� �                                    ?� �                                     �  x                                     �  p                                    � �                                    � �                                     �  p                                     �  `                                    �  �                                    �  �                                     �  `                                     �  @                                    �@ �                                    �@ �                                     �  @                                                                             �� �                                    �� �                                                                                                                      �   �                                    �   �                                                                                                                       �                                         �                                                                                                                           t                                         t                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      