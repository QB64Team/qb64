��d  |J� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         ����������������������������������������������������������������������������������������������������������������������������������������������������������������������� �                                       ������������������������������������������������������������������������������������������������������������������������������ ����������������������������������������������������������������������������������������������������������������������������������������������������������������������� �������������������������������������������                                       o���������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                  �  p ������������������������������������������������������������������������������������������������������������������������������    �      �   �    >          ���� p �������������?������������������� ����������������������������          ��p ����������������?����������������������������   ��     �   �   ��         ��� �p ������ ���������?���� ?����������0� �������������������������           ����������� ���������?�������������������������   �     `  �  ���          � �p ����������������?���  ������������� ������������������������            ���������������������?�������������������������   <�     p`  �  ��     ;+ � ��� �p �������������������   ��������i��� �����������������������       ;+ � �������������������������     ;+ � ��������   �      ��  �  ��     $��T �����p �����������������  ��������������������������������������       $��T �p ����������������������     $��T ��������  �~     �      ��     $��T ����p �����?�������?������    ������WR���������������������������?        $��T �p �������?�������?������?��     $��T ��������  ��A�� �   ���    $��T ����p ���������?���w���    �����W^����������������������������        $��T �p �����������?���w�������    $��T ��������  �����  x�>   ���    $��T ����p �����??��x?��������  ?������������������������������������             �p �������??��x?�����������    $��T ��������   � :9���  ���   ��    $��� ����p ��������ps?����� �      $��� �����������������������������               ����������ps?���������    $��� ���������   ?�bq�� ���              ����p ��������p�?���f1��� �          ������������������������������              ����������p�?���f1�����          ���������   ��a�9� ;�             �    � p ������9�a�����<����         �  ������������������������������              ���������9�a�����<�������       �  ���������    ���7  3�                      p �������>c������x�����              ���������������������������������������������������>c������x���������������������������  ���8~ 8w                      p ������<ǁ���ǈ�������               ��������������������������������������������������<ǁ���ǈ����������������������������  ��0x 0�8                      p �������|χ������������              ���������������������������������������������������|χ��������������������������������  > >�0� a�p                      p ��������y�=������������������������������������������������������������������������������y�=�������������������������������  p ��`� ��8�                      p ������	�q�9���<3������������������������������������������������������������������������	�q�9���<3���������������������������  `�1�`� 8��1�                      p ������9�c�1���13������������������������������������������������������������������������9�c�1���13���������������������������  ����� ���3�                      p ������?��'������������������������������������������������������������������������?��'���������������������������  ���@p �y�`                      p ������?�����w������������������������������������������������������������������������?�����w���������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p ����������    ������     ������    �����������������������������������������������������������������������������������������                                      p �����������������������������������������������������������������������������������������������������������������������������                                      p �����������������������������������������������������������������������������������������������������������������������������                                      p �����������������������������������������������������������������������������������������������������������������������������                                      p �����������������������������������������������������������������������������������������������������������������������������                                      p �����������������������������������������������������������������������������������������������������������������������������   "r�       ����      ' �<        p �����ݍ�|�������c|�������������_��������ݍ�|��������c|�������������������������ݍ�|��������c|����������������������   "��       ����      /��>        p �������|��������A|���>��_�����ϟ����������|��������A|��������_������������������|��������A|��������_�������������   "��       ����      /��>        p �������|��������A|�������_�����������������|��������A|��������_������������������|��������A|��������_�������������   "��     p ����     /��>       p �������|�������A|�������_�����~�����������|��������A|��������_������������������|��������A|��������_�������������   "�     � ��     " (��       p ������u�������w�]}���������_�����|����������u�������w��]}����������_�����������������u�������w��]}����������_�������������   >�      ��      蠀       p ������u����������]}��������_����������������u����������]}���������_�����������������u����������]}���������_�������������   >�      ���x     ��       p ������u����������]|?�������_����������������u����������]|?��������_�����������������u����������]|?��������_�������������   >�      ����     ��       p ������u���������]|?������_����������������u����������]|?�������_�����������������u����������]|?�������_�������������   >�       ����     ��    	   p ������u�������߿�]|?������_����������������u����������]|?�������_�����������������u����������]|?�������_�������������   "�     @ �� �     (��    �  p ������u������￿�]}��������_������{���������u����������]}���������_����������������u����������]}���������_������������   "�     � �� �    " (��       p ������u��������]}��������_�����~����������u���������]}���������_�����������������u���������]}���������_�������������   "��     � ����     /��>       p ������~������A�������A�����~����������~�������A��������A�����������������~�������A��������A�������������   "��       ����      /��>        p ������~��������A�������A����������������~��������A��������A�����������������~��������A��������A�������������   "��       ����      /��>        p ������~��������A���>��A�����ϟ���������~��������A��������A�����������������~��������A��������A�������������   "s�       ����      '>�<        p �����݌~�������c�������������_��������݌~��������c�������������������������݌~��������c����������������������                                      p �����������������������������������������������������������������������������������������������������������������������������                                      p �����������������������������������������������������������������������������������������������������������������������������                                      p �����������������������������������������������������������������������������������������������������������������������������                                      p �����������������������������������������������������������������������������������������������������������������������������                                      p �����������������������������������������������������������������������������������������������������������������������������                                      p ����������    ������     ������    �����������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p ����                                 �����������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p ����������    ������     ������    �����������������������������������������������������������������������������������������                                      p �����������������������������������������������������������������������������������������������������������������������������                                      p �����������������������������������������������������������������������������������������������������������������������������                                      p �����������������������������������������������������������������������������������������������������������������������������                                      p �����������������������������������������������������������������������������������������������������������������������������                                      p �����������������������������������������������������������������������������������������������������������������������������   "r�@      ����      ' �        p �����ݍ�}�������c|�������������_��������ݍ�}��������c|�������������������������ݍ�}��������c|����������������������   "��@      ����      /��>        p �������}��������A|���>��_�����ϟ����������}��������A|��������_������������������}��������A|��������_�������������   "��@      ����      /��>        p �������}��������A|�������_�����������������}��������A|��������_������������������}��������A|��������_�������������   "��@     ����     /��>       p �������}�������A|�������_�����x�����������}��������A|��������_������������������}��������A|��������_�������������   "�@    0 �� �     (��     �  p ������u���������]}��������_�����ww���������u����������]}���������_����������������u����������]}���������_������������   >��    0 �� �     蠀      �  p ������u������Ͽ�]}�������_������{���������u���������]}��������_����������������u���������]}��������_������������   >��    P ����     ��<     �  p ������u�����ﯿ�]|?������_������{���������u���������]|?�������_����������������u���������]|?�������_������������   >��    P ����     ��>       p ������u�����ﯿ�]|?������_����������������u���������]|?�������_�����������������u���������]|?�������_�������������   >��    � ����    $ ��>       p ������u������o��]|?������_����������������u������o��]|?�������_�����������������u������o��]|?�������_�������������   "��    � ��     > (��"       p ������u��������]}���������_����������������u��������]}����������_�����������������u��������]}����������_�������������   "� @     ��      (��"       p ������u���������]}���������_�����w����������u����������]}����������_�����������������u����������]}����������_�������������   "��@     ����     /��>    �  p �������������A�������A�����pw�����������������A��������A������������������������A��������A������������   "��@      ����      /��>        p ��������������A�������A������������������������A��������A�������������������������A��������A�������������   "��@      ����      /��>        p ��������������A���>��A�����ϟ�����������������A��������A�������������������������A��������A�������������   "s�@      ����      '>�        p �����݌�������c�������������_��������݌��������c�������������������������݌��������c����������������������                                      p �����������������������������������������������������������������������������������������������������������������������������                                      p �����������������������������������������������������������������������������������������������������������������������������                                      p �����������������������������������������������������������������������������������������������������������������������������                                      p �����������������������������������������������������������������������������������������������������������������������������                                      p �����������������������������������������������������������������������������������������������������������������������������                                      p ����������    ������     ������    �����������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p ����                                 �����������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p ����������    ������     ������    �����������������������������������������������������������������������������������������                                      p �����������������������������������������������������������������������������������������������������������������������������                                      p �����������������������������������������������������������������������������������������������������������������������������                                      p �����������������������������������������������������������������������������������������������������������������������������                                      p �����������������������������������������������������������������������������������������������������������������������������                                      p �����������������������������������������������������������������������������������������������������������������������������   "r��      ���p      ' �        p �����ݍ�|������c|��������������_��������ݍ�|�������c|��������������������������ݍ�|�������c|�����������������������   "���      ����      /��>        p �������|�������A|���>��_�����ϟ����������|�������A|��������_������������������|�������A|��������_�������������   "���      ����      /��>        p �������|�������A|�������_�����������������|�������A|��������_������������������|�������A|��������_�������������   "���    p ����     /��>       p �������|������A|�������_�����x�����������|�������A|��������_������������������|�������A|��������_�������������   "�      � �� �    " (��"    �  p ������u�������w�]}�w�������_�����ww���������u�������w��]}�w��������_����������������u�������w��]}�w��������_������������   >�       �� �     蠀"     �  p ������u����������]}�w������_������{���������u����������]}�w�������_����������������u����������]}�w�������_������������   >� @     ����     ��>     �  p ������u����������]|?������_������{���������u����������]|?�������_����������������u����������]|?�������_������������   >� @    0 ���p     ��>       p ������u�������Ͽ�]|?�������_����������������u����������]|?��������_�����������������u����������]|?��������_�������������   >� @     ����     ��     �  p ������u����������]|?������_������{���������u����������]|?�������_����������������u����������]|?�������_������������   "� @     �� �     (��     �  p ������u����������]}�w�������_������{���������u����������]}�w��������_����������������u����������]}�w��������_������������   "� �    � �� �    " (��    �  p ������u��}����w�]}�w�������_�����ww���������u������w��]}�w��������_����������������u������w��]}�w��������_������������   "�    p ����     /��>       p ������}������A�������A�����x�����������������A��������A������������������������A��������A�������������   "�      ����      /��>        p ������}�������A�������A�����������������������A��������A������������������������A��������A�������������   "�      ����      /��>        p ������}�������A���>��A�����ϟ����������������A��������A������������������������A��������A�������������   "s      ���p      '>�<        p �����݌}������c��������������_��������݌�������c��������������������������݌�������c�����������������������                                      p �����������������������������������������������������������������������������������������������������������������������������                                      p �����������������������������������������������������������������������������������������������������������������������������                                      p �����������������������������������������������������������������������������������������������������������������������������                                      p �����������������������������������������������������������������������������������������������������������������������������                                      p �����������������������������������������������������������������������������������������������������������������������������                                      p ����������    ������     ������    �����������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p ����                                 �����������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p ���������������������                �����������������������������������������������������������������������������������������                                      p ������������������������������������������������������������������������������������������������������������������������������                                      p ������������������������������������������������������������������������������������������������������������������������������                                      p ������������������������������������������������������������������������������������������������������������������������������                                      p ������������������������������������������������������������������������������������������������������������������������������                                      p �����������������������������������>_�����������������������������������������������������������������������������������������      �   � �                       p ������������?�������������������������������������������������������������������������������?�����������������������������      �  � ?�                       p �����������?������������������������������������������������������������������������������?�����������������������������        � �                       p ��������������������������������������������������������������������������������������������������������������������������         ��0                   �  p ��������������?�������������������w���������������������������������������������������������?��������������������������           �                  @  p �������������������������������������������������������������������������������������������������������������������������          �                   @  p �������������������������������������������������������������������������������������������������������������������������      �! � ��c�               @  p �����������=����<9�����������������������������������������������������������������������=����<9�����������������������      �g�� ����               #�  p ����������~9���8���������������{������������������������������������������������������~9���8����������������������       [�  ?�Lg��               D@  p ��������������x��f�������������ﻻ�����������������������������������������������������������x��f�����������������������      `��  ��n3                �@  p �����������3���3'�����������������{����������������������������������������{����������������3���3'������������������{�������      @�1� ��0l&`              @  p �����������3��?'ϓٟ������������������������������������������������������������������������3��?'ϓٟ�����������������������      �1�c� ��0�|`              �  p ��������?�9�w��?�#����������������w���������������������������������������������������?�9�w��?�#�����������������������      �1�Ø ��`��                    p ��������?�s<g���'����������������������������������������������������������������������?�s<g���'������������������������     �c���da��                    p ���������rp��?�O9�����������������������������������������������������������������������rp��?�O9������������������������     �c��>fg0�                    p ����������d������s������������������������������������������������������������������������d������s������������������������      ��0��~~`��                   p ���������9��� �����������������>_������������������������������������������������������9��� ��������������������������      �0�0  8<`�                   p ���������9������ß����������������������������������������������������������������������9������ß�����������������������                                      p ������������������������������������������������������������������������������������������������������������������������������                                      p ������������������������������������������������������������������������������������������������������������������������������                                      p ������������������������������������������������������������������������������������������������������������������������������                                      p ���������������������                �����������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������         �      0                   p ������������������������������������������������������������������������������������������������������������������������������               0     �            p ������������������������������������������������������������������������������������������������������������������������������               0     �            p ������������������������������������������������������������������������������������������������������������������������������         �8�<��6<l�<���g�         p ������������������������������������������������������a��'�Ó���$��������������������������������������������������������         �3m���<fl�3f훶l�         p �����������������������������������������������������̒O�'Ù��g̙dI�?�������������������������������������������������������         ?0�>��8~l�0f͛6o�         p ��������������������������������������������������������?�3'ǁ��gϙ2dɐ?�������������������������������������������������������         0`f��<`l�0f͛6l          p �������������������������������������������������������矙3'ß��gϙ2dɓ��������������������������������������������������������         3m�f�p6f8�3f͛6��         p ������������������������������������������������������̒O�3�ə��g̙2d�?�������������������������������������������������������         8�>�`3<0�<��3�`        p ���������������������������������������������������������3�������3$�d�������������������������������������������������������                `  0                  p �������������������������������������������������������������������������������������������������������������������������������               �  �                  p �����������������������������������������������������������?������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p ���������������������������������������������������������������������������������������������������������������������������������������������������������������������� ��                                      ?����������������������������������������������������������������������������������������������������������������������������� ����������������������������������������������������������������������������������������������������������������������������������������������������������������������� �������������������������������������������                                       ��������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         ������������������������������������������������������������������������������������������������������������������������������