�'k  �0� }                                                                                                                                                                                                          8                                                                                                                           `                                                                         �                                               �                                                ��                                              ��                                               �x                       �                      �`                                               ��                        `                      ��                                               ��                                             ��                                               ���                                             ���                                              ��x                       �                     ��`                                              ���                        `                     ���                                              ���                                            ���                                              '����                                           &���                                             y��x                      �                    y��`                                             ~� �                       `                    |� �                                             | �                    �                      }| �                                             � ��                    @                      � ��                                            � �x                    @  �                   � �`                                            �  �                        `                   ^  �                                             �  �                                           ^  �                                             o  ��                                          /  ��                                            o  �x                      �                   /  �`                                            7�  �                       `                   �  �                                            7�  �                                         �  �                                            �  ��                                         �  ��                                           �  �x                      �                  �  �`                                           ������                       `                  �  ��                                           ������                                        ������                                           �  ���                 ���                   �  ���                                          ������x                      �                 ������`                                          ������                  �     `                 ������                                          ������                 �                      ������                                          ��������                 @                       �������                                          �    �x                 @     �                 �    �@                                          �     �                        `                 ^     �                                          �     �                                        ^     �                                          o     ��                                       /     �                                          o     �x                     �                /     ~@                                         7�    ��                      `                �    ?�                                         7�    �                     �                �    ?�                                         �    w��                     �                �     7��                                        �    ��x                     @�               �    �`                                        �    ���                     @ `               �     ߘ                                        �     ���                                     �     ���                                        �     ����                                     �     ����                                       �     m��x                    @�              �     E�`                                       x     m��               �     @ `              x     E�                                       x     7`�              �     �               x      �                                       �     7`��              @     �                �       ��                                      �     ��x              @       �              �     @�`                                       �     � �                       `              ^     @ �                                       �     � �                                    ^     � �                                       o     � ��                                    /     � ��                                      o        �x                      �             /        �`                                      7�        �                       `             �        �                                      7�        �                                   �        �                                      �        ��                                   �        ��                                     �        �x                      �            �        �`                                     �         �                       `            �         �                                     �         �                                  �         �                                     �         ��                                  �         ��                                    �         �x                      �           �         �`                                    x          �            �           `           x          �                                    x          �           �                      x          �                                    �          ��           @                       �          ��                                   �          �x           @           �           �          �`                                    �           �                        `           ^           �                                    �           �                                  ^           �                                    o           ��                                  /           �                                   o           ��                                  /           ��                                   7�           �                                  �           ?�                                   7�           ��                                �           ?�                                   �           ��                                �           ?�                                  �           �x                      �         �           ?�`                                  �           ���                       `         �           ?�                                  �           ���                               �           _��                                  �           ����                               �           o���                                 �          ���x                      �        �           ��`                                 x          � �         �              `        x           � �                                 x          � �        �                      x           � �                                 �          � ��        @                       �          � ��                                �          � �x        @              �        �          � �`                                 �          �  �                        `        ^          �  �                                 �          �  �                               ^          �  �                                 o          �  ��                              /          �  ��                                o          �  �x                      �       /          �  �`                                7�         �   �                       `       �         �   �                                7�         �   �                             �              �                                �         `   ��                �           �          @   ��                               �            �x                �    �      �              �`                               �              �                `     `      �         �    �                               �         #�    �               �           �         @    �                               �         #�    �                �     �     �         @    �                               �         #�    ��               �            �         @                                   x               ��      �         `           x         �     �                             x              ��      �         �     �     x                �                       �     �         `     ��      @         �     �      �               �                       �     �         �    ��      @                �      �                �                       �      �         �    ?��                              F         �    �                              �         �   ���                                       �    8                                         �   ���                      8        3         �   ǀ                                         �   ~?�                      �        1         �   ?�                                �        �  ���                                �        �   q��                                �        �  ��                       p          �        �  ��                                 �        �  ��                      �         @        �  �                                 �        � ���                                         �  ���                                 �        � ?�                       �          .�        � �                                  �        ����                                 .�        � 8��                                  �        ����                      8           .�        ����                                  �    ����~?�                    �           Q       �|?�                                   ��   ?��������                                 N�    �� �q��                                   ?��   ?� ����                      p             ;�   ?� ���                                    �������������             |   |                 ��       ��                                     ?�����������             �                       ?����������                                     �|   |  ��              ��������               �|   |  �~               |   |                  �����������                                      ����������p                                      �����������                                      �����������                                       ?���������                |   |                   ?��������|                                        ���������                |   |                   ���������                                        ��   �                  ����                   �    �                                           �������                        �                  ������@                                           ~    �                        @                  ~    �                                                 �                                                 �                                                 `                                                 `                                   