�h  �z��                 `                                              `                                              `                                              `                                             �` 0                                           �` 0                                           �` 0                                           �` 0                                            ` 0                                            ` 0                                            ` 0                                            ` 0                                           g�8<��ny����<��<                               g�8<��ny����<��<                               g�8<��ny����<��<                               g�8<��ny����<��<                               3lٰf��l��m���f                               3lٰf��l��m���f                               3lٰf��l��m���f                               3lٰf��l��m���f                               �o�0f�������0>͛~                               �o�0f�������0>͛~                               �o�0f�������0>͛~                               �o�0f�������0>͛~                                                                                                                                       �l03f�����͛0f͛`                                                                                                                                                                                           �lٰ3f́�l͛m�0f͛f                                                                                                                                                                                           g�<���fy���0>��<�                                                                                                                                                                                                                                                                                                                                                                                                                           �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ?��                ��                ��                                                                                                                                                                       � |                �               | �                                                                                                                                                                      x  �             �                �  <                                                                                                                                                                     �   8                 �             8   �                                                                                                                                                                                     0                 �    `                                                                                                                                                                    0    �            �                                                                                                                                                                                         �     `                �                                                                                                                                                                                                          `           0     �                                                                                                                                                                                   0                 �      `                                                                                                                                                                                   @                                                                                                                                                                                                 �          �                                                                                                                                                                                         �       `                �                                                                                                                                                                                                          @                                                                                                                                                                                                                             �                                                                                                                                                                                                  @        @                                                                                                                                                                                                   �                                                                                                                                                                                          @                                                                                                                                                                                                   �        �                                                                                                                                                                                         @         @                                                                                                                                                                                                 �                           �                                                                                                                                                                                                         @                                                                                                                                                                                                                           �                                                                                                                                                                                                          �                                                                                                                                                                                              @          @                                                                                                                                                                                              �                                                                                                                                                                                      @                                                                                                                                                                                                      @                                                                                                                                                                                                 �      �                                                                                                                                                                                                �      �                                                                                                                                                                                    @           @                                                                                                                                                                                       @     @           @                                                                                                                                     @                                                   �     �                             �                                                                                                                    �            @                  @                        �                             �                                                                             @                  @                               @                  �                                                    @                                                                             @                  �                               �                  �                                                    @                                                                             �                  �                               �                                                                                         �                                                            �                                                                                                                                          �                                                                                                                                                                                                       �                                                                                                                                                  @                                       @            @                                                                                                @                                                 �                                       @            @                                                                                                �                                                                                        @            @                                                                                                                                                                                        @            @                                                                                                                                                                                          �                                                                                                                                                                                                       �                                                                                                                        �                                               �                �          �     �             �                                   �                              �                               `                                   �           �                �          �                   �                                   �            `                 �                  �            P                                   �           �                �          �                  �                                  �             H                 �                 �             �                                  �           <          @     �               p           �                 8                 �            �                 �                 �            �                                  @                     @     �               �           �                 |                 �             �                 �                              �                                  .�           s�         @     7�               1�           ��                o                 ?�            �                 /�                 @            O�                ?                 ]<           ��         @     /��              c�           ��                0��                            #                                  �            �                `�                �           �<         @     _��              ���          ��                q��                ���           P�                .                 9            
��                 �               t?�          ��         @     ��<             ���          ��                a��               �?�           L0                �p�                r�            <�                @��               ���          ���        @     ���             �<          |��               ���               ���           �                |0                �0�           ??�              ���               ���          ���        @    ���            ??�          ?�              ����              ���           ��                �               �0           ��               ��?�              ���          3��<        @    ���            ���         ���              ��?�              ����          - 0�              � �               �           *��              ���              O�?�         7�?�        @    ���<            ����         >���              ���              ��?�          	 0              � 0�                �           ��              �3�              .����         g����       @    ��?�            1���<         =���             �3�              ?����          Z �              �0              @0�          T<?�              ��              3�3�         ����       @    ����           #��?�         }�?�             ���             ?�3�          �  �              �               � 0          1� ��             `?�             =��         �� �<       @    ����           ߀��        {� ��             ?`?�             ����         �  0�             �� �              "           �� 3�             ` ��             ��?�        �� ?�       @    �� �<           ���        �� 3�             ` ��             ��?�         %  0             �� 0�               �          a� �              � 3�             !� ��        x ��      @    �� ?�           �� �<        w� ��             o� 3�             >� ��         h�              �@ 0             $�  0�         1� ?�            7� �             @ހ 3�        x ��           �� ��      �     �� ?�         � ?�             �� ��             �� 3�         (�  �             @              @	  0         "�  ��            K� ?�            �/@ �        �  �<            N� ��      �     ;� ��        �  ��             O� ?�             ?@ ��         H  0�               �             ��          @�  3�            �  ��            @ ?�       �  ?�            �  �<      �     � ��        �  3�             �  ��             @ ?�        @H  0               0�            �  �         @z  �            �  3�            �  ��        �  ��           x  ?�      �     �  �<         �  ��            �  3�             �  ��        @$               �  0            @  0�        �z  ?�            �  �            �  3�        �  ��           x  ��     �     �  ?�         �  ?�            �  ��            �  3�        �$   �              �              @  0        �=   ��             �  ?�           �  �        o   �<          �  ��     @     �  ��@       }   ��            �  ?�            �  ��       �   0�             H   �                       =   3�           @ �   ��           �  ?�       o   ?�          �   �<     @     �  ��@       }   3�            �   ��            �  ?�          0           @ H   0�               �        �  �           � z   3�            �   ��       7�  ��           �   ?�     @     x   �<@       >�  ��            �   3�            �   ��       	              � $   0             �   0�       �  ?�          � z   �          @ �   3�       7�  ��           �   ��     @     x   ?�@       >�  ?�            �   ��           �   3�       	    �           � $             @  �   0       @  ���           =  �?�         �  �  ��       �����8           o������           ������       �����            }����?�           ������       �   0�               �          �  H          ���3�           =��� ��           ����?       ������           o�����            �������       ���3�            }��� ��           ����?       �  ?�0              �0�           H  ��       �����           �����           ��� O          ��           4   ��            �  ���       �����            ?�����            ���� O       �����            �����            /�����       ����            �����           ���        ������           7������           ������        ����             ?�����            ����           ��              ?�                ��       ���� @           ����            ?���        ������           ������           o�����        ���� @            ����             ���           ��              ?��              ��       �                                 8       �     ������           ������           o�����        �                                   x            �����           �����            �����       ������           �����             �����  �     �����           ������           7�����        ������            �����             ?�����        �                                               �                 �             @   �      @     x    @           �               7�           �                 �                 >�             �                 @             @   	              �                 �             �   @      @     �    @           �               �           �                 �                 @             H                               �   �          @  �              @  �                @            �    �      �     �               �           �                 �                 @          @  H              @                   �          @  z              �  �                �             �    �      �     x               �            �                 �                 �          @  $              �   �                @          �  z              �  �                �            �          @     x               �            �                 �                 �          �  $              �   �                @          �  =                 �                �            o          @     �               �            }                 �                 �          �                   H                             =                 �                �            o                �          �     �             }                 �                 �                             H                             �                z                 �            7�               �          @     x   @         >�                 �                 �            	                 $                  �            �                z            @    �            7�               �                 x   �         >�                 �                 �            	                 $            @     �            @                =            �     �            �               o                 �   �         @                 }                 �            �                            �     H            @                =                 �            �               o   @            �            @                 }                 �            �                                 H            �                �                z       �     �                7�  �             �            �                 >�                 �            @                	                 $            �                 �                 z       @     �  @             7�               �            �                 >�                 �            @                 	                  $            �                 @                 =             �  �        �     �               o            �                 @                 }                              �                             �            @    @                 =            �          @     �               o            �                 @                 }                         @    �                             �            �    �                 �           x                �          �     7�            �                 �                 >�            �            �    @                 	             �            �    �                 �           x               �          @     7� @          �                 �                 >�             �            �    @                 	              �                �                 @           �               �                 � �          �                 �                 @             H                                  �        @    �                �                 @           �               � @              �           �                 �                 @        @    H                                  �        @    z                 �                 �       �     � `              x�              �            �                 �                 �        @    $                  �                 @        �    z                 �                 �             � �          �    x               �            �                 �                 �        �    $                  �                 @        �    =                  �                 �            o           @    �               �            }                 �                 �        �                      H                              =                  �                 �            o           0    �           �    �`            }                 �                 �                              H                               �                 z                 �            7�                �`           0    y�            >�                 �                 �             	                  $                  �             �                 z                 �        �    7�                ߀               ~             >�                 �                 �             	                  $                  �                               8                  �        0    �            �    n                �                               x                 �                                                 @                                                  �                         0    x             �   �                               `                 �                                                                                                                �   8                 �             8   �                                                                                                                                                                     x  �             �                �  <                                                                                                                                                                      � |                �               | �                                                                                                                                                                       ?��                ��                ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      � `�  ��         ̀`             �         0                                                                                                                                                              0    ��         l `�             0     0                                                                                                                                                                 0    ��          `�             0     0                                                                                                                                                                 1�n�><��;`<��<     �|�y�<��y�      ��͹��3π                                                                                                                                                            1��lٻ�����f     ͳv�Ͷf���      ͳ3m�m�7m�n�                                                                                                                                                            1��lٳ>����>͛~      m�f���~��͘      3?m��3�f6l�                                                                                                                                                            1��lٳf����f͛`      m�f���`�f͘      30m�3c6l�                                                                                                                                                            1��lٳf���`f͛f     m�f�ͶfͶ͘      �3m�m�6m�l�                                                                                                                                                            1��f�3>��30>��<     ͟f`y�<��y�      �m�͙�g3��                                                                                                                                                                                                                                                                                                                                                                                      �        >                                                                                 