��g  @  ���>��00��>  ��@@��  ����  ���  �    ���   �� � ���G��6��?������?�������>��  �����        ���>��00��>"�"����EDED����ğ��"�2������  @��   �� � ���G��6��?������?�������>��  �����        ���>��00��>  ��AED���FG�Gď������������PP���
��#����h.�<���2r���8<|x���>�?�������>��  �����        ���>��00����  ����@@����@@�������������������� ����� ����@ ���� @����  ���� 0 ����� ����                ��  �     P�P'�'�� K�[��@��_�@TT_�@��_�@$4_�@/�  P�      �� �                        ��  �     �   $H� @H$�@ O�@ O�@ O�@ $O�@ H'�  �       �� �                ���������>�>�>�>���������������������������������������������>�>�>�>��������          ��  ����  O� �>  >�   �  `
@�  @ �@ @ �@ @ �@ @ �@ @ �  `
 �   �> >��� O�  ��  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      