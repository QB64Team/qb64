��d   ��!                                                                 ?������������������                                    ?������������������                                                                                           ?������������������                                    @                                                      @                                                      ?������������������                                    ������������������                                    �                                                      �                                                      ������������������                                    �������������������                                                                                                                                                �������������������                                   �                 �                                   �����������������                                    �����������������                                    �                 �                                   �                 �                                   ?�����������������                                    ?�����������������                                    �                 �                                   �                 �                                   �����������������                                    �����������������                                    �                 �                                   @                 �                                   ������������������                                    ������������������                                    @                 �                                   �                 �                                   !?�����������������                                    !?�����������������                                    �                 �                                   =�                 �                                   B?�����������������                                    B                                                     =��m�$�I#m��rI$�6�l�                                   {�                 �                                   ������������������                                    �@                                                    {����   ����   ���                                   �                  �                                  ������������������                                   �                                                    ����   ����   ���                                  �                  �                                  ����������������������������������                                   ����������������                  �6�m�$�I#m��rI$�6�l�                                  �                  �����������������                  #������������������                                 "                                                  ����   ����   �������������������                  �                  �����������������                  G������������������                                 D                                                  ����   ����   �������������������                  p                  �����������������                  �������������������                                 �                                                  r6�m�$�I#m��rI$�6�l�����������������                  �                  �                                 !�����������������������������������                 !                 �����������������                 ����   ����   ���                                 =�                  �               �                 B?����������������������������������@                 B                  ����������������@                 =����   ����   ���               �                 {�               �  �               �                 �����������������������������������                  �@               | ����������������                  {�6�m�$�I#m��rI$���l�               �                 �               W� �               �                �����������������������������������                �              � ����������������                 � ���   ����  ����               �                �               � �                �                ����������������T�����������������                               ������������������                � ���   ����  ����                �                �               |` �                x                #����������������)?������������������                "               ��                �                ܒ6�m�$�I#m��rI$���l�$�I#m��rI$�6�m� x                �               �` �                <                G����������������������������������                D               U�                �                � ���   ����  ����   ����   ��� <                p               �� �                                �������������������������������������                �               U`                �                p ���   ����  ����   ����   ���                 �               �� �                                !���������������檏�������������������               !               Up                ��               �6�m�$�I#m��rI$���l�$�I#m��rI$�6�m�$                =�               �� �                �               B?����������������������������������@               B                Up                 �@               =� ���   ����  ����   ����   ��� �               {�               U� �                �               ����������������� �������������������                �@               Up                 |                {� ���   ����  U���   ����   ��� �               �                U` �                �              ����������������� ?������������������              �               UP                 >               �$�6�m�$�I#m��rI$�U{l�$�I#m��rI$�6�m�$��              �                U  �                 �              ����������������� ?������������������                              UP                               �  ���   ����  U��   ����   ���  �              �                Up �                 x              #����������������� �������������������              "                U`                 �              �  ���   ����  U��   ����   ���  x              �                T@ �                 <              G����������������� ?�������������������              D                U`                 �              ��m�$�H�m�ܒI$���mUd���m�ܒI$���m�$�H�h<              p                ` �                               ������������������ ?�������������������              �                U@                 �              w���  ����   ���U` �����   ����  ��              �                � �                               !����������������� ��������������������             !                U�                 ��             ����  ����   ���U� �����   ����  ��              =�                ր �                 �             B?�������������������������������������@             B                 �                   �@             =��m�$�H�m�ܒI$���oפ���m�ܒI$���m�$�H�m�             {�                 |  �                 �             ��������������������������������������              �@                 �                   |              {����  ����   ����  �����   ����  ����             �                     �                 �            ���������������������������������������            �                                     >             ����  ����   ����  �����   ����  ����            �                     �                  �            ���������������������������������������                                                             ��m�$�H�m�ܒI$���m�$���m�ܒI$���m�$�H�m��            �                     �                  x            #����������������������������������������            "                                     �            �����  ����   ����  �����   ����  ���x            �                     �                  <            G����������������������������������������            D                                     �            �����  ����   ����  �����   ����  ���<            p                     �                              �����������������������������������������            �                                      �            u��m�$�H�m�ܒI$���m�$���m�ܒI$���m�$�H�m�            �                     �                              !�����������������������������������������           !                                      ��           �����  ����   ����  �����   ����  ���            =�                     �                  �           B?����������������������������������������@           B                                        �@           =�����  ����   ����  �����   ����  ����           {�                     �                  �           �����������������������������������������            �@                                       |            {���m�$�H�m�ܒI$���m�$���m�ܒI$���m�$�H�m���           �                      �                  �          �����������������������������������������          �                                      >           �����  ����   ����  �����   ����  �����          �                      �                   �          �����������������������������������������                                                           �����  ����   ����  �����   ����  �����          �                      �                   x          #������������������������������������������          "                                        �          ܍��m�$�H�m�ܒI$���m�$���m�ܒI$���m�$�H�m��x          �                      �                   <          G������������������������������������������          D                                        �          �����  ����   ����  �����   ����  ����<          p                      �                             �������������������������������������������          �                                        �          p����  ����   ����  �����   ����  ����          �                   �  �                             !�������������������������������������������         !                   |                    ��         䍶�m�$�H�m�ܒI$���m�$���m�ܒI$���m�$�H�m��          =�                  W� �                   �         B?������������������������������������������@         B                   �                     �@         =�����  ����   ����� �����   ����  �����         {�                  � �                   �         ��������������������T���������������������          �@                  ��                    |          {�����  ����   ����� �����   ����  �����         �                   |` �                   �        ��������������������)?���������������������        �                  ��                    >         �$���m�$�H�m�ܒI$���o����m�ܒI$���m�$�H�m�܁�        �                   �` �                    �        �����������������������������������������                           U�                            � ����  ����   ����� �����   ����  ���� �        �                   �� �                    x        #��������������������������������������������        "                   U`                    �        � ����  ����   ����� �����   ����  ���� x        �                   �� �                    <        G�������������������檏����������������������        D                   Up                    �        �$���m�$�H�m�ܒI$��������m�ܒI$���m�$�H�m�ܐ<        p                   �� �                            �������������������������������������������        �                   Up                    �        p ����  ����   ����� �����   ����  ����         �                   U� �                            !�������������������� ������������������������       !                   Up                    ��       � ����  ����   ���U� �����   ����  ����         =�                   U` �                    �       B?�������������������� ?����������������������@       B                    UP                     �@       =�$���m�$�H�m�ܒI$���Ut���m�ܒI$���m�$�H�m�ܒ�       {�                   U  �                    �       ��������������������� ?����������������������        �@                   UP                     |        {� ����  ����   ���Up �����   ����  ���� �       �                    Up �                    �      ��������������������� ����������������������      �                   U`                     >       �  ����  ����   ���Up �����   ����  ���� �      �                    T@ �                     �      ��������������������� ?����������������������                          U`                           ��rI$�6�m�$�I#m��rI$�U{l�$�I#m��rI$�6�m�$�I#m��      �                    ` �                     x      #��������������������� ?�����������������������      "                    U@                     �      ����   ���   ����  U��   ����   ���   ��x      �                    � �                     <      G��������������������� �����������������������      D                    U�                     �      ����   ���   ����  U���   ����   ���   ��<      p                    ր �                           ����������������������������������������������      �                    �                      �      u��rI$�6�m�$�I#m��rI$���l�$�I#m��rI$�6�m�$�I#m�      �                     |  �                           !����������������������������������������������     !                     �                      ��     ����   ���   ����   ����   ����   ���   ��      =�                        �                     �     B?����������������������������������������������@     B                                              �@     =����   ���   ����   ���   ����   ���   ���     {�                        �                     �     �����������������������������������������������      �@                                            |      {���rI$�6�m�$�I#m��rI$�6�l�$�I#m��rI$�6�m�$�I#m���     �                         �                     �    �����������������������������������������������    �                                            >     ����   ���   ����   ���   ����   ���   ����    �                         �                      �    �����������������������������������������������                                                     �����   ���   ����   ���   ����   ���   ����    �                         �                      x    #������������������������������������������������    "                                              �    �m��rI$�6�m�$�I#m��rI$�6�l�$�I#m��rI$�6�m�$�I#m��x    �                         �                      <    G������������������������������������������������    D                                              �    �����   ���   ����   ���   ����   ���   ���<    p                         �                          �������������������������������������������������    �                                              �    w����   ���   ����   ���   ����   ���   ���    �                         �                          !�������������������������������������������������   !                                              ��   �m��rI$�6�m�$�I#m��rI$�6�l�$�I#m��rI$�6�m�$�I#m��    =�                         �                      �   B?������������������������������������������������@   B                                               �@   =�����   ���   ����   ���   ����   ���   ����   {�                         �                      �   �������������������������������������������������    �@                                              |    {�����   ���   ����   ���   ����   ���   �����   �                          �                      �  �������������������������������������������������  �                                               >   �#m��rI$�6�m�$�I#m��rI$�6�l�$�I#m��rI$�6�m�$�I#m��A�  �                          �                       �  �������������������������������������������������                                                    �����   ���   ����   ���   ����   ���   �����  �                          �                       x  #��������������������������������������������������  "                                                �  �����   ���   ����   ���   ����   ���   ����x  �                       �  �                       <  G��������������������������������������������������  D                       |                        �  �#m��rI$�6�m�$�I#m��rI$���l�$�I#m��rI$�6�m�$�I#m��p<  p                      W� �                         ���������������������������������������������������  �                      �                        �  p����   ���   ����  ����   ����   ���   ����  �                      � �                         !�����������������������T�������������������������� !                      ��                       �� �����   ���   ����  ����   ����   ���   ����  =�                      |` �                       � B?�����������������������)?�������������������������@ B                       ��                        �@ =�#m��rI$�6�m�$�I#m��rI$���l�$�I#m��rI$�6�m�$�I#m��r� {�                      �` �                       � �������������������������������������������������  �@                      U�                        |  {�����   ���   ����  ����   ����   ���   ����� w                       �� �                       � ���������������������������������������������������� ��                      U`                        > w ����   ���   ����  ����   ����   ���   ����� v                       �� �                        � ������������������������檏������������������������� �                       Up                         vI#m��rI$�6�m�$�I#m��rI$���l�$�I#m��rI$�6�m�$�I#m��r@� t                       �� �                        x ��������������������������������������������������� �                       Up                        � t ����   ���   ����  ����   ����   ���   ���� x p                       U� �                        < ������������������������� ��������������������������� �                       Up                        � p ����   ���   ����  U���   ����   ���   ���� < p                       U` �                         ������������������������� ?�������������������������� �                       UP                        � rI#m��rI$�6�m�$�I#m��rI$�U{l�$�I#m��rI$�6�m�$�I#m��rH p                       U  �                         ������������������������� ?����������������������������                       UP                        ��p ����   ���   ����  U��   ����   ���   ����  p                       Up �                        �������������������������� ��������������������������@�                       U`                         �@p ����   ���   ����  U��   ����   ���   ���� �p                       T@ �                        �������������������������� ?�������������������������� �                       U`                         | u�ܒI$���m�$�H�m�ܒI$���mUd���m�ܒI$���m�$�H�m�ܒI$����p                       ` �                        �������������������������� ?���������������������������                       U@                         >w��   ����  ����   ���U` �����   ����  ����   ���p                       � �                         �������������������������� ���������������������������                       U�                         w��   ����  ����   ���U� �����   ����  ����   ���p                       ր �                         x������������������������������������������������������                       �                          �u�ܒI$���m�$�H�m�ܒI$���oפ���m�ܒI$���m�$�H�m�ܒI$���xp                        |  �                         <����������������������������������������������������                        �                          �w��   ����  ����   ����  �����   ����  ����   ��<p                           �                         ������������������������������������������������������                                                   �w��   ����  ����   ����  �����   ����  ����   ��p                           �                         ������������������������������������������������������                                                  �u�ܒI$���m�$�H�m�ܒI$���m�$���m�ܒI$���m�$�H�m�ܒI$���p                           �                         ������������������������������������������������������                                                   �w��   ����  ����   ����  �����   ����  ����   ��p                           �                         ������������������������������������������������������                                                   bw��   ����  ����   ����  �����   ����  ����   ���p                           �                         ������������������������������������������������������                                                    "u�ܒI$���m�$�H�m�ܒI$���m�$���m�ܒI$���m�$�H�m�ܒI$���\p                           �                         ������������������������������������������������������                                                    "w��   ����  ����   ����  �����   ����  ����   ���p                           �                         ������������������������������������������������������                                                    "w��   ����  ����   ����  �����   ����  ����   ���p                           �                         ������������������������������������������������������                                                    "u�ܒI$���m�$�H�m�ܒI$���m�$���m�ܒI$���m�$�H�m�ܒI$���\p                           �                         ������������������������������������������������������                                                   "w��   ����  ����   ����  �����   ����  ����   ���p                           �                         ������������������������������������������������������              ������������                         "w��   ����  ��            �����   ����  ����   ���p              �������������                         ����������������            ��������������������������                                                     "u�ܒI$���m�$�H�_��������������m�ܒI$���m�$�H�m�ܒI$���\p              ?�������������                         ����������������            ��������������������������              @                                      "w��   ����  �������������������   ����  ����   ���p              �������������                         ����������������            ��������������������������              �                                      "w��   ����  ������������������   ����  ����   ���p              �                                      ������������������������������������������������������             �������������                         "u�ܒI$���m�$�H��            �m�ܒI$���m�$�H�m�ܒI$���\p             �                                      ������������������������������������������������������             �������������                         "w��   ����  ��            ����   ����  ����   ���p             �                                      ���������������?���������������������������������������             ?�������������                         "w��   ����  ��            ����   ����  ����   ���p             �                                      ���������������_���������������������������������������             _�������������                         "u�ܒI$���m�$�Hנ            �m�ܒI$���m�$�H�m�ܒI$���\p             `                                      ������������������������������������������������������             ��������������                         "w��   ����  �`            ����   ����  ����   ���p             �                                      ������������������������������������������������������             !�������������                         "w��   ����  ��            ����   ����  ����   ���p             =�                                      ������������������������������������������������������             B�������������                         "u�ܒI$���m�$�H��            �m�ܒI$���m�$�H�m�ܒI$���\p             {�                                      ������������������������������������������������������             ��������������                         "w��   ����  {�            ����   ����  ����   ���p             ��                                      �����������������������������������������������������            ������������������������              "w��   ����   ��                       �  ����   ���p            ��            �����������              ���������������������������          ���������������            �������������                        "u�ܒI$���m�$�I��            ������������$�H�m�ܒI$���\p            ��            �����������              �������������� �������������          ���������������             �������������                        "w��   ����  ��            ������������  ����   ���p            ��            �����������              ��������������@�������������          ���������������            @�������������                        "w��   ����  ��            ������������  ����   ���p            �                                     ������������������������������������������������������            �������������������������              "rI#m��rI$�6�m��                       6�m�$�I#m��rI$�p            ��                                     �������������� ���������������������������������������            ! �������������������������             "p ����   �����                       ���   ����  p            =��                       �             �������������� ��������������������������������������            B ������������������������@             "p ����   �����                       ����   ����  p            {��                       �             �������������� ������������������������?��������������            � ������������������������              "rI#m��rI$�6�m{��                       ��m�$�I#m��rI$�p            ���                       �             ������������� ��������������������������������������            ������������������������             "p ����   �����                       ����   ����  p            ���                        �             ������������� ��������������������������������������            ������������������������             "p ����   �����                        ����   ����  p            ���                        x             ������������� ���������������������������������������            �������������������������             "rI#m��rI$�6�l���                        z�m�$�I#m��rI$�p            ���                        <             ������������� ���������������������������������������            �������������������������             "p ����   �����                        =���   ����  p            ���                                     ������������� ?���������������������������������������            ?�������������������������             "p ����   �����                        ���   ����  p            ���                                     �������������                         ���������������                                    ��            "rI#m��rI$�6�l���                        [m�$�I#m��rI$�p            ���                        �            ������������� @                       ��������������            @                       �@            "p ����   �����                        ���   ����  p            ��                         �            ������������� �                       �?�������������            �                       �             "p ����   ����                         ���   ����  p            ��                         �            �������������                        ��������������                                   �            "rI#m��rI$�6�l��                         �m�$�I#m��rI$�p            ��                          �            �������������                         ��������������                                    �            "p ����   ����                          ���   ����  p            ��                          x            �������������                         ��������������                                    �            "p ����   ����                          {��   ����  p            ��                          <            �������������                         ?��������������                                    ?�            "rI#m��rI$�6�l��                          =m�$�I#m��rI$�p            ��                                      �������������                         ��������������                                    �            "p ����   ����                          ��   ����  p            ��                                      �������������                          ��������������                                     �            "p ����   ����                          ��   ����  p            �                                      �������������@                         ��������������           @                         �            "rI#m��rI$�6�l�                          m�$�I#m��rI$�p            �              �                       ��������������                         ��������������           �             �          �            "p ����   ���                           ��   ����  p            �              �                       �������������                          ��������������                         �          �            "p ����   ���                           ��   ����  p            �              �                       �������������                        ��������������                         �           �            "rI#m��rI$�6�l�                        m�$�I#m��rI$�p            �              �                       �������������            �           q�������������                         �           q            "p ����   ���            �           ��   ����  p            �           �  �                       �������������            @A           1�������������                      �  �           1            "p ����   ���            @A           ��   ����  p            �          �  �                       �������������            `@           �������������                     �  �                       "rI#m��rI$�6�l�            `@           m�$�I#m��rI$�p            x          �  �                       ��������������            `8@           �������������           �          �  �                       "p ����   ��x            `8@           ��   ����  p            <          � ��                       ��������������            p(�8           �������������           �          � ��                       "p ����   ��<            p(�8           ��   ����  p                      ��                         ��������������           @p8�8           �������������           �          ��                         "rI#m��rI$�6�l           Pp8�8           m�$�I#m��rI$�p                      � �  >                      ���������������         �x0�8@          �������������           ��         � �  >                      "p ����   ��          �x0�8@          ��   ����  p            �         ��^                       ��������������@           xp�9�          �������������            �@         ��^                       "p ����   ���          p��9�          ��   ����  p            �         ���\ ��                     ��������������            x`��          �������������            |          ���\ ��                     "u�ܒI$���m�$��           ����          �H�m�ܒI$���\p            �         �� ���                     ��������������         x`��          �������������            >         �� ,��                     "w��   ����  �         �`�           ����   ���p             �         � ���                     ��������������          �a��$          �������������                     �   ��                     "w��   ����   �         �`�,           ����   ���p             x          �  ���                     ���������������          ����          �������������            �          �   ��                     "u�ܒI$���m�$�@x          ���          �H�m�ܒI$���\p             <          @  ��                     ���������������         ����� >         �������������            �          @  ��                     "w��   ����   <         �����>          ����   ���p                       @� ��                     ���������������         ߸py0�"         �������������            �          @� ��                     "w��   ����            ��py0�"          ����   ���p                        � >��                     ����������������        _�rg!�           !�������������            ��          �  ��         !            "u�ܒI$���m�$�H         _�pg!�           �H�m�ܒI$���\p             �          � >          <            ���������������@       �Fpb��           C�������������             �@          �           C            "w��   ����  �       �Fpb��           < ����   ���p             �            >?�         z            ���������������        �Cx�F�           ��������������             |             ?�         �            "w��   ����  ��       �Cx�f��         z ����   ���p             �       � 8  �         �            ���������������        C��t�n         	�������������             >       �    �        	            "u�ܒI$���m�$�H��        C��t�o�         ��H�m�ܒI$���\p              �       � |   �        �            ���������������        ?��x��         �������������                    �     �                    "w��   ����  ��        ?��x���        � ����   ���p              x       � �    �        �            ����������������        ?��h�8         #�������������             �       �     �        "            "w��   ����  �x       ?�h�8�        � ����   ���p              <       À�   x        �            ����������������        ����?`         G�������������             �       � (   x        D            "u�ܒI$���m�$�H�<       })��?`x        ��H�m�ܒI$���\p                     ���   >8        p            ����������������        ���I��         ��������������             �       �    >8        �            "w��   ����  �       ?�I��8        p ����   ���p                     �|            �            �����������������       ���G��        !�������������             ��                    !            "w��   ����  �       ?��G��        � ����   ���p              �       �8           =�            ����������������@      ?����_��        B?�������������              �@             w        B             "u�ܒI$���m�$�H��      ?���_��        =ĒH�m�ܒI$���\p              �      8�            {�            ����������������        ������        ��������������              |       8              �@            "w��   ����  ���      8������        {� ����   ���p              �      p    � >        �             ����������������       �������       ��������������              >      p      >       �            "w��   ����  ���      p������        �  ����   ���p               �      p   �        �             ����������������       ������       ��������������                    p                          "u�ܒI$���m�$�H�`�      p�����       �$�H�m�ܒI$���\p               x      �   ��  �      �             �����������������      ������       #��������������              �      �   �@  �      "             "w��   ����  ��x      ����N]���      �  ����   ���p               <      �  ��  C�      �             �����������������      �����        G��������������              �      �  �   C�      D             "w��   ����  ��<      ��� ��      �  ����   ���p                    � ��  ��      p             �����������������      �5�@��@       ���������������              �     � 
�   ��      �             "u�ܒI$���m�$�H�l     ��1�@�A�      q$�H�m�ܒI$���\p                    � �  A�      �             ������������������      �?t����        !��������������              ��    �  �   A�      !             "w��   ����  ��     �� t�����      �  ����   ���p               �    � ?�� ��      =�             �����������������@      ?tG����       B?��������������               �@    �  ��   �      B              "w��   ����  ���    �? tG����      =�  ����   ���p               �    ��?�� ��      {�             �����������������       >?�����       ���������������               |     ���  �      �@             "u�ܒI$���m�$�H�m��    �>v��?��      {�$�H�m�ܒI$���\p               �       ?�� � �      �              �����������������    ��;����      ���������������               >       
 �   �     �             "w��   ����  ����    ��w�?��      �   ����   ���p                �    � ?�  � �     �              �����������������    �w/���      ���������������                   � $�    �                   "w��   ����  ����    ��w/�?��     �  ����   ���p                x    �    � `     �              ������������������    �?�?�����     #���������������               �    �        `     "              "u�ܒI$���m�$�H�m�x    �� �?����     ��$�H�m�ܒI$���\p                <    �   @  `     �              ������������������    �%�?��� �     G���������������               �    � 
      `     D              "w��   ����  ���<    ��!�?��� �     ��  ����   ���p                    �    ��  p     p              ������������������    '�'�� �     ����������������               �    �    �  `     �              "w��   ����  ���    �'�'� �     w�  ����   ���p                    �@   ]�  �     �              �������������������    �����     !���������������               ��   �@   �  �     !              "rI#m��rI$�6�m�$�H    �������     �6�m�$�I#m��rI$�p                �   ��   �  �     =�              ������������������@    ��t8     B?���������������                �@   ��   �  �     B               "p ����   ���   �   ���t8�     =����   ����  p                �   �@  �  �     {�              ������������������    ���� @     ����������������                |    �@   �  �     �@              "p ����   ���   �   ����� B�     {����   ����  p                �   � � �� �     �               ������������������   ������     ����������������                >   �    �� �    �              "rI#m��rI$�6�m�$�I�   ������ �     �6�m�$�I#m��rI$�p                 �   � � ���    �               ������������������   ����� x     ����������������                   �    ���                   "p ����   ���    �   ���?��px�    � ���   ����  p                 x   � �����    �               �������������������   ?����     #����������������                �   �   ���    "               "p ����   ���    x   �?�>�t�    � ���   ����  x                 <   ������    �               �������������������    q����      G����������������                �   �   ���    D               "zI#m��rI$�6�m�$�I <   �q�<�p�    ��6�m�$�I#m��rI$�<                    ���/���    p               �������������������    �?����     ������������������                �   �  ����    �               "< ����   ���      ��0|����    p ���   ����                      ��w� �    �               ��������������������   ��t� �     !�����������������                ��   � @� �    !               " ����   ���      ��x�Ԉ ��    � ���   ����                   �  � �#� �    =�               �������������������@  ������    B?������������������                �@   �  �� �    B                "I#m��rI$�6�m�$�I#�  ��������    =Ē6�m�$�I#m��rI$��               �  �   �     {�               ������������������   ��� ���    ������������������@               |    p   � �    �@               "�����   ���   ��  ��� ����    {� ���   ����  �            �   �  �     �     �                �?�����������������  � �� ��@   ������������������            �   >   p     � �   �               "�����   ����  ��  � �� ��G�    �  ���   ����  �            @    �  �          �                �����������������  �@�� ��     ������������������           �      8       �                   "�#m��rI$�6�m��I#`�  �@�� �� �   �$�6�m�$�I#m��rI$� �                 x  �       8   �                �������������?�����  �@�� ��  8   #������������������           �   �   8       �   "                " �����   ����  �x  �@�� �� �   �  ���   ����   x                <  �     @ <8   �                �������������������  �@w ��� 8   G�������������������           �   �          ?�   D                " x����   ����  �<  �@w ���?�   �  ���   ����   <                x  �       88   p                �������������������  �@s��� 8   ��������������������           ?�   �          ?�   �                " =#m��rI$�6�m���I#lx  �@s���?�   q$�6�m�$�I#m��rI$�                 �  �      x0   �                ������������������  �@p8��� 0   !�������������������           �            �   !                " ����   ����  ��  �@p8����   �  ���   ����                  �  ��     �p   =�                <������������������  �  `$��p p   B?��������������������          ��      �     ��   B                 B ����   ����  ��  �� `$��p��   =�  ���   ����  < �              �  �� ?�  �p   {�                x������������ ����2  �  @$�0 p   ��������������������@         ��   2   � ?�  ��   �@                � �m��rI$�6�m���I#k�  �� @$�0��   {�$�6�m�$�I#m��rI$x �            �  �  �� ?�  �p   �                 ���?����������  ����b  �  D$�0  p  �������������������          ���  b   � ?�  ��  �                �����   ����� ��  �� D$�0��   �   ���   ����  � �            @  <  �� ?�  ��  �                �������������  ����  �  @ X0  �  �������������������         ���  �    � ?�  �                    �����   ����� �<  �� @ X0��  �   ���   ���� �  �               |  ��     �  �                �������������  ?���  �� @ P0  �  #�����������������2��         ���  !�    |    �   "                2  �m��rI$�6�o���I#^|  �� @ P0��  �I$�6�m�$�I#m��rI#�  x              <�  ��    | �  �                ��������������  ���  �� ` D   �  G�����������������b���         ���  C        �   D                b  {����   ����� ��  �� ` D ��  �   ���   ���� �  <              y�  ���   ��  p                <�������������  ���  �� @ H  �  ����������������������         ?���  �    ?�   ��   �                �  =����   ����� y�  ���@ H!���  p   ���   ���� <           �    ��  ���   ��  �                |������������π ?��  ��   p  �  !��������������������         p��     �   ��   !                !�  m��rI$�6����I"��  ���  p#���  �I$�6�m�$�I#m��rI|           0` @ ��  ���   ��  =�                <��������������` ��  ��   `  �  B?���������������������        ϟ��     �   ��   B                 C  ���   ����� ��  ���  `���  =�   ���   ���� <�  �        @ � ��   ��� � �  {�                y������������@ ���0   ��      �  ���������������������@       ���  0    �� ���   �@                �  ����   ����� ��   ���� ����  {�   ���   ���� y�  �        �  ��   ��� ��  =                 �����?�������� ���`   ��     �  ���������������������        ���  `    �� ���                    Ͷ�rI$�6�����I'��   ���� ����  =rI$�6�m�$�I#m��rH��  �        �  ?�   ���� ?���                  ������������ ����   ���    ��  ��������������������       ���  �     � ?��   �                  ����   ����  ?�   ���� ?����  �   ���   ������   �         �   �������                   ��?�������������   ��   �   ������������������0 ?��       ���  !�    �����   ��               0    ����   ����  �   ��������   `   ���   ������   x        �  <��   �x?��    �               �����������������    �x       �����������������`@���       �{�  C     �������   �@               `@   zI$���m�?���m����   ��������   ���m�$�H�m�ܒI$����   <        �  y��   ?�� � >   �               ? ���������������    ?�� � >   �?���������������������       ?�{�  �     �?����   �                ��   <  ����?�����y��   ?��������   �����  ����   �?            �   ���   �� � |   �               ~ ������������?��    �� � |   ����������������� ���       �{�       �����   �               !�      ������������   ��������   �����  ����   �~            @ ���   ��?��  �    �               <� �������������    ��?��  �   ����������������� ����      ����       � ��    �               C    I$���m�����m����   ��������    ���m�$�H�m�ܒI$���    �        � ���   ���� �    x               y� ��������� ����0    ���� �   ������������������ ���@     ���  0      ?� ��    ��               �    � �������������   ��������    {����  ����   y�    �        	  ���   ��    �    <               ��  ���?������ �	���`    ��    �   �����������������  ���      ���  `      �����    ��                  � �������������   ��������    =����  ����   ��    �          ?��   ��    �                  ��  �������� @����    ��    �   ����������������  ��     ���  �      �����    �                  �$���m�����m�?��   ��������    ��m�$�H�m�ܒI$���     �        d  ��   ��    �                  ��  ?�������� 0���    ��    �   ?����������������0   ?��     ���  !�      �����    ?��             0      � ������������   ��������    ���  ����   ��     x       �  <���   ��    �    �             ��  ��������� ���     ��    �   ���������������`@  ���     ���  C        �����    �@             `@     x �������������   ��������    ����  ����   ��     <          y���    ���   ��    �   �        ?   ���������  ���       ���   ��   �?���������������  ���     ?���  �         ���     �    �        ��     =$���m�����my���    ��������    ��m�'�H�m�ܒI$�?                 ��߀    ��  �     �   �        ~   ���������  ?��  @    ��  �    ���������������   ���     ���   @      ���     �   �        !�       �����������߀    ������     ���������   ~              @ ���     ��  ?�      �   �        <�   ��������   �� P�    ��  ?�    ��������������   ����    ���  P�      ���     �   �        C       �����������     ������      ���������   <�      �       � ��v     �����      x   �        y�   ��������  ���0 �     �����    ���������������   ���@    ?��  0 �        �      ��   �        �      ����m�����k��v     ������      z�m�?�H�m�ܒI$y�      �        ���     ������      <   
        ��    ���?����� ���`     ������     ��������������    ���     ��  `                 ��   ;�             ������������     ������      =���?�����   ��      �        ?��     ������         ;�       ��    ������� ����     ������     ��������������    ��    ��  �                 �   4             ���������?��     ������      ���?�����  ��       �        ��      ������         >>       ��    ?������� ���      ������     ?��������������0     ?��    ��  !�                 ?��  0       0        ��m���H�^��      ������      [m�?�H�m�ܒI#��       x        <���      ?����       �  <
       ��    �������� ���  �     ?����      ������������`@    ���    ��  C  �                �@  0       `@       x�����������      ?����       ���>����  ��       <        y����     ����       �  8       ?     �������� ���  @     ����      �?�������������    ���    ��  �  @                �   0       ��       <�������y����     ����       ���<����  ?                 �����     ����       �         ~     �������� ?��         ����      ������������     ���     ��                     �         !�        ���m���H������     ����       �m�<H�m�ܒI~              @ �����      ?��         �  8       <�     �������� �� @       ?��       ����#��������     ����    �  @                 �         C        �����������      ?��         ���<����  <�        �     � ����      ��         x  �       y�     �����������0 �       ��       �������������     ���@    ?  0 �                 ��  �       �        �����?������      ��         {�������  y�        �      �����                  <  �       ��      ���?��������`                   ������������      ���       `                   ��  �              Ͷ�m��Hן����                  =m�'�H�m�ܒH��        �      ?����                            ��      �����������                   ������������      ��      �                   �                  ����� �?����                  ��  ���� ��         �      ����                            ��      ?����������                   ?������������0       ?��       !�                   ?��         0          ����� �����                  �  ���� ��         x       <�����                  �         ��      �����������   
                 �����������`@      ���       C   
                 �@         `@         y��m�$�H������                  ��$�H�m�ܒG��         <       y�����                  �         ?       �����������                    �?������������      ���       �                    �          ��         =����  y�����                  ߀  ���� ?                 ������                  �         ~       ����������    "                 �����������       ���          "                 �         !�          ����   ������                  �  ���� ~                ������                   �         <�       ���������� @  B                 �����������       ����      @  B                 �         C          6�m�$�I������                   ��$�H�m�ܒ<�          �     ����|                   x         y�       ���������0 �  �                 ������������       ���@     0 �  �                 ��         �          ����  ����|                   {�  ���� y�          �     ������                   <         ��        ���?������`                    �����������        ���      `                    ��                  ����  ������                   =�  ���� ��          �     ?�����                           ��        ���������                    ����������        ��     �                    �                  �$�6�m�?�����                   6�m�$�I#m��           �     �����                           ��        ?��������                    ?����������0         ?��     !�                    ?��       0            �  ��������                   ���   ���           x     <������                   �       ��        ���������                     ���������`@        ���     C                     �@       `@           x  ���������                   ����   ���           <     y������                   �       ?         ���������                     �?����������        ���     �                     �        ��           =$�6�my������                   ��m�$�I#o?                 �������                   �       ~         ��������                        ���������         ���                            �       !�              ���������                   ����   �~                �������                    �       <�         �������� @  @@                  ���������         ����    @  @@                  �       C              ���������                    ����   ��            �   ����                     x       y�         �������0 �  ��                  ����������         ���@   0 �  ��                  ��       �            ��6�k����                     z�m�$�I#y�            �   ������                     <       ��          ���?����`                      ���������          ���    `                      ��                  � ��������                     =���   ��            �   ?�����                           ��          �������                      ��������          ��   �                      �                  � ��?�����                     ���   ��             �   �����                           ��          ?������                      ?��������0           ?��   !�                      ?��     0              ��6�^�����                     [m�$�I#��             x   <������                     �     ��          �������                       �������`@          ���   C                       �@     `@             x ��������                     ���   ��             <   y������                     �     ?           �������                       �?��������          ���   �                       �      ��             < �y������                     ���   ?                 �������                     �     ~           ������                          �������           ���                            �     !�              �6��������                     �m�$�I~                �������                      �     <�           ������ @  @@                    �������           ����  @  @@                    �     C               ��������                      ���   <�              � ����                       x     y�           �����0 �  ��                    ��������           ���@ 0 �  ��                    ��     �              ������                       {��   y�              � ������                       <     ��            ���?��`                        �������            ���  `                        ��                  �6ן�����                       =m�$�H��              � ?�����                           ��            �����                        ������            �� �                        �                  ��?�����                       ��  ��               � �����                           ��            ?����                        ?������0             ?�� !�                        ?��   0                �������                       �  ��               x <������                       �   ��            �����                         �����`@            ��� C                         �@   `@               z6�������                       ��$�G��               < y������                       �   ?             �����                         �?������            ��� �                         �    ��               <y������                       ��  ?                 �������                       �   ~             ����                            �����             ���                            �   !�                ~�������                       ��  ~                �������                        �   <�             ���� @  @@                      �����             ���� @  @@                      �   C                5�������                        ��$�<�                �����                         x   y�             ���|0 �  ��                      ������             ���D0 �  ��                      ��   �                �����                         {�  y�                ǟ�����                         <   ��              ���8`                          �����              ���(`                          ��                  ן�����                         =�  ��                �?�����                           ��              ���                          ����              ���                          �                  �?�����                         �$���                 ������                           ��              ?���                          ?����0               ?���                          ?�� 0                  ������                         ~ ��                 |������                         � ��              ���                           ���`@              ���                           �@ `@                 |������                         � ��                 9������                         � ?               ���                           �?����              ���                           �  ��                 9������                         �$�?                  ������                         � ~               ���                             ���               ���                             � !�                  ������                         � ~                  ������                          � <�               ���   @@                        ���               ���   @@                        � C                  ������                          � <�                  ���                           x y�               ��� � ��                        ����               ��� � ��                        �� �                  ���                           x�y�                  ��?��                           < ��                ��� �                          ���                ��� �                          ��                  ��?��                           =���                  ����                           ��                �� �                          ��                �� �                          �                  ����                           ���                  ����                           ��                ?�� �                          ?��0                 ?�� �                          ?��0                   ����                           [��                  ����                           ���                �� �                          �x`@                �� �                          �H`@                  ����                           ���                  ����                           �?                 �� '�                          �0��                �� '�                          �0��                  ����                           �?                   ����                           �~                 �� C�                            ��                 �� C�                            ��                   ����                           �~                   �  ��                            ��                 �� ��@@                          �                 �� ��@@                          �                   �  ��                            ��                   �                               y�                 �� ���                          ��                 �� ���                          ��                   �                               y�                   �  ~                             3�                  �� �                            ��                  �� �                            ��                   �  ~                             3�                   �  |                             �                  � ?�                            �                  � ?�                            �                   �  |                             �                   �  x                             �                  ?� �                            ?�                   ?� �                            ?�                    �  x                             �                   �  p                             �                  � �                            �@                  � �                            �@                   �  p                             �                   �  `                                                �  �                            ��                  �  �                            ��                   �  `                                                 �  @                                                �@ �                            �                   �@ �                            �                    �  @                                                                                                     �� �                            �                   �� �                            �                                                                                                                             �   �                            �                   �   �                            �                                                                                                                              �                                 �                    �                                 �                                                                                                                               t                                 p                    t                                 p                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                