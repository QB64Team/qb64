�l  �z��                 `                                              `                                              `                                              `                                             �` 0                                           �` 0                                           �` 0                                           �` 0                                            ` 0                                            ` 0                                            ` 0                                            ` 0                                           g�8<��ny����<��<                               g�8<��ny����<��<                               g�8<��ny����<��<                               g�8<��ny����<��<                               3lٰf��l��m���f                               3lٰf��l��m���f                               3lٰf��l��m���f                               3lٰf��l��m���f                               �o�0f�������0>͛~                               �o�0f�������0>͛~                               �o�0f�������0>͛~                               �o�0f�������0>͛~                                                                                                                                       �l03f�����͛0f͛`                                                                                                                                                                                           �lٰ3f́�l͛m�0f͛f                                                                                                                                                                                           g�<���fy���0>��<�                                                                                                                                                                                                                                                                                                                                                                                                                           �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ?��                ��                ��                                                                                                                                                                       � |                �               | �                                                                                                                                                                      x  �             �                �  <                                                                                                                                                                     �   8                 �             8   �                                                                                                                                                                                     0                 �    `                                                                                                                                                                    0    �            �                                                                                                                                                                                         �     `                �                                                                                                                                                                                                          `           0     �                                                                                                                                                                                   0                 �      `                                                                                                                                                                                   @                                                                                                                                                                                                 �          �                                                                                                                                                                                         �       `                �                                                                                                                                                                                                          @                                                                                                                                                                                                                             �                                                                                                                                                                                                  @        @                                                                                                                                                                                                   �                                                                                                                                                                                          @                                                                                                                                                                                                   �        �                                                                                                                                                                                         @         @                                                                                                                                                                                                 �                           �                                                                                                                                                                                                          @                                                                                                                                                                                                                             �                                                                                                                                                                                                           �                                                                                                                                                                                              @          @                                                                                                                                   @                                                           �                                                                                           @                                                  �                                         @                                                                                                           �                                                  �                                         @                                                                                                           �                                                                                      �      �                                                                                                                                                                                                �      �                                                                                                                                                                                    @           @                                                                                                                                                                                     @     @           @                                                                                                                                   @                                                 �     �                             �                                                                                                                  �                                                       �                             �                                                                                                                                                                                                      @                                                                                                                               @                                                                       @                                                                             @                                                  @                                                                                          �                                                            @                                                  �                  @                                                                       �                                                            �                  @                               �                  �                                                                        �                                                            �                  �                                                  �                  @                                       @            @                                                                              �                  @                                                 �                                       @            @                                                                                                �                                                                                        @            @                                                                                                                                                                                        @            @                                                                                                                                                                                         �                                                                                                                                           �                                                           �                                       �                                                                                 h                  �                  �                             @          �                    @                  0                  �                                                              l                 x                 �                             �          �      `             D                 8                                                                                   �                 ~                                               �          �      �             �                 x                                                                                   �                 �                 8                       @                     �            �                  �                                                                                 �                 �                 x            @          @                     �                            �                 0                                                                �                 �                 �            @          @                                                  	�                 `                                                                �                �                 1�            �          @                                 (                 �                  �                                                                �                ��                c��           �          @                                 /�                �                 A�                                                                �?�               7���               ǃ�          �         @                    8|           X>                '��                ��                                                               ���               /��              ���          >         @      �              p�          _��               ?�              �                                                               ���              _��?�             ���          �        @       �             �           ��               N�<              ���                                                              ����              �����             ?���                  @        <            �  �         ����              ����             ��                                                              ����             ����?�            ���           �       @     @  �           �           w��              <���<             7���                                                             ����            �����            ����                 @     �   <              �        p���            9���À            g��                                                             7����           ���~            �����           �      @     �   �                     "���            y���p             ׀���                                                            7� ���           �� ?���           �� ��?       @         @        p             �       "� ��            �� ?��            �� ��8                                                            o�  ��~           �� ���           �� ���      @   �     @                       8       E�  ��p            �� ���           � ��                                                           �  ���           �x  ?�?           #�  ���           p     @      �   �                     ^  ��            �x  ?�8           �  ���                                                           ^   ���           �x  ���          @�  �                        �    8     �          �       ^   ���           Ix  ��            �  �                         �                 @              o   �<          �   ��          ��  ���          �            @         �                  /   �0           �   ��           �  ��                                          �               o   ��          �   �0          �   ?��           2            @     �     �                  /   ��            �   �0           �   ?��                                                         7�   �           �   ��          x   �                              8     �      �     �       �   �            ^   ��           x   �                                                         @7�   �           �    ?�          x    ��                                  �      �             �   �            ^    ?�           x    ��      @                                                 @�   �           o    �          �    �                                @      @     @       �   �            /    �            �    �      @                                                 ��    8           o     �          �    �                                @      @     @       �    8            /     �            �    �      �                                                 ��               7�                 �     �                                @            @       �                �                 ^     �      �                                                  �                 7�              @  �                                      @            @       �                 �                 ^                                               @               �                 �              �  o                                                   �       �                 �                 /                                               �               �               @ �                o                                                   �       �                 �                 /                             @                                x               � �                7�            �                                      �       x                 �                 �                            �                                x               � �                7�            �                    @                       x                 �                 �                            �                                �                �                �            @                    @                        �                 �                 �                                                            �                �                �      �      @                     �                        �                 �                 �                                                             �                x                 �      �                        �    �                        ^                 x                 �                                                              �                x             @   �      @           @            �                            ^                 x                 �                                            @                 o                �             �   �      @          @            @                            /                  �                 �                                            �                  o                �                �                 �      �      @                            /                  �                 �                                                               7�                �                x                 �      �                       �            �                 ^                 x                                                            @  7�                 �                x                      @                       �            �                 ^                 x          @                                                  @  �                 o                �                      @                      @            �                 /                  �          @                                                  �  �             @   o                �                                       �      @             �                 /                  �          �                 @                                �  �             �   7�                 �                                      @          @         �                 �                 ^          �                 �                                   �             �   7�           @     �                                                  �         �                 �                 ^                           �                @                  �                �           �     o                                                 �         �                 �                 /                                           �                  �                �                o                               @                         �                 �                 /                                                             x                �                7�      �      �                   �                         x                 �                 �                                                            x                �                 7�      @      �  @                                         x                 �                 �                                                             �                �                 �             @  �        �                                  �                 �                 �                                                             �                �                 �            @          @                                  �                 �                 �                                                              �                x                 �                              �          �                   ^                 x                 �                                                              �                 x                 �                             �          @       @           ^                 x                 �                                                               o                 �                 �                            @                   �           /                  �                 �                                                                o            @    �                 �                            @ @                           /                  �                 �                          @                                      7�           �     �                 x       �      `                �               �            �                 ^                 x                          �                                 @    7�                 �                 x              �          �                      �            �                 ^                 x        @                                                   @    �                 o                 �                       @                     @            �                 /                  �        @                                                   �    �                 o                 �                       0                �     @`            �                 /                  �        �                                                   �    �                 7�                 �                            `           0     !�            �                 �                 ^        �                                                        �                 6                  �        �    `                	�                &             �                                   X                                                                                                     `        0    �            �                                                                                                                                                                                                        0                 �    `                                                                                                                                                                    �   8                 �             8   �                                                                                                                                                                     x  �             �                �  <                                                                                                                                                                      � |                �               | �                                                                                                                                                                       ?��                ��                ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      � `�  ��         ̀`             �         0                                                                                                                                                              0    ��         l `�             0     0                                                                                                                                                                 0    ��          `�             0     0                                                                                                                                                                 1�n�><��;`<��<     �|�y�<��y�      ��͹��3π                                                                                                                                                            1��lٻ�����f     ͳv�Ͷf���      ͳ3m�m�7m�n�                                                                                                                                                            1��lٳ>����>͛~      m�f���~��͘      3?m��3�f6l�                                                                                                                                                            1��lٳf����f͛`      m�f���`�f͘      30m�3c6l�                                                                                                                                                            1��lٳf���`f͛f     m�f�ͶfͶ͘      �3m�m�6m�l�                                                                                                                                                            1��f�3>��30>��<     ͟f`y�<��y�      �m�͙�g3��                                                                                                                                                                                                                                                                                                                                                                                      �        >                                                                                 