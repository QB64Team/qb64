��b   ˀ� ��                 ��������������������������������������� @                �                    �                                                                                                                      @                                                                              @                  ��                 ��������������������������������������� @                �                    �                                                                                                                      @                                                                              @                  ��                 ��������������������������������������� @                �                    �                                                                                                                      @                                                                              @                  ��                 ��������������������������������������� @                �                    �                                                                                                                      @                                                                              @                  ��                 ��������������������������������������� @                �                    �                                                                                                                      @                                                                              @                  ��                 ��������������������������������������� @                �                    �                                                                                                                      @                                                                              @                  ��                 ��������������������������������������� @                �                    �                                                                                                                      @                                                                              @                  ��                 ��������������������������������������� @                �                    �                                                                                                                      @                                                                              @                  ��                 ��������������������������������������� @                �                    �                                                                                                                      @                                                                              @                  ��                 ��������������������������������������� @                �                    �                                                                                                                      @                                                                              @                  ��                 ��������������������������������������� @                �                    �                                                                                                                      @                                                                              @                  ��                 ��������������������������������������� @                �                    �                                                                                                                      @                                                                              @                  ��                 ��������������������������������������� @                �                    �                                                                                                                      @                                                                              @                  ��                 ��������������������������������������� @                �                    �                                                                                                                      @                                                                              @                  ��                 ��������������������������������������� @                �                    �                                                                                                                      @                                                                              @                  ��                 ��������������������������������������� @                �                    �                                                                                                                      @                                                                              @                  ��                 ��������������������������������������� @                �                    �                                                                                                                      @                                                                              @                  ��                 ��������������������������������������� @                �                    �                                                                                                                      @                                                                              @                  ��                 ��������������������������������������� @                �                    �                                                                                                                      @                                                                              @                  ��                 ��������������������������������������� @                �                    �                                                                                                                      @                                                                              @                  ��                 ��������������������������������������� @                �                    �                                                                                                                      @                                                                              @                  ��                 ��������������������������������������� @                �                    �                                                                                                                      @                                                                              @                  ��                 ��������������������������������������� @                �                    �                                                                                                                      @                                                                              @                  ��                 ��������������������������������������� @                �                    �                                                                                                                      @                                                                              @                  ��                 ���������������������������������������� @                �                                                                                                   ���������������������������������������� @                                                                              @                  ��                                                          @                �                                                                                                                                            @                                                                              @                  ��                                                          @                �                                                                                                                                            @                                                                              @                  ��                                                          @                �                                                                                                                                            @                                                                              @                  ��                                                          @                �                                                                                                                                            @                                                                              @                  ��                                                          @                �                                                                                                                                            @                                                                              @                  ��                                                          @                �                                                                                                                                            @                                                                              @                  ��                                                          @                �                                                                                                                                            @                                                                              @                  ��                                                                            �                                                            @                                                                              @                                                                              @                  ��                                                                            �                                                            @                                                                              @                                                                              @                  ��                                                                            �                  �������������������������������������������                                    �������������������������������������������                                    �������������������������������������������                  ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            �                                                                                                                                                                                                                                                ��                                                                            � �����������������������������������������������������������������������������                                                                                                                                                                 ��������������������������������������������������������������������������������                                                                                                                                                              p                                                                                ��������������������������������������������������������������������������������                                                                              p                                                                              �                                                                                ��������������������������������������������������������������������������������                                                                              �*�                                                                            T                                                                                ��������������������������������������������������������������������������������                                                                              �$�                                                                            $                                                                                ��������������������������������������������������������������������������������                                                                              �(�                                                                            D                                                                                ��������������������������������������������������������������������������������                                                                              p                                                                              �                                                                                ��������������������������������������������������������������������������������                                                                                                                                                              p                                                                                ��������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            