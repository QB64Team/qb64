��]  |J� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         ����������������������������������������������������������������������������������������������������������������������������������������������������������������������� �                                       ������������������������������������������������������������������������������������������������������������������������������ ����������������������������������������������������������������������������������������������������������������������������������������������������������������������� �������������������������������������������                                       o���������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������         �       �                 p ������������������?���������������������������������������������������������������������������������?������������������������        �       � � �             p ������������������?�������������������������������������������������������������������������������?����������������������        `      �   0     0        p ���������������������������������������������������������������������������������������������������������������������������        `          `     `        p �����������������������������������������������������������������������������������������������������������������������������        0@      �   �     �        p ����������Ͽ������������������������������������������������������������������������������Ͽ�����������������������������        `       �  ��     �        p ����������������������� �����?�������������������������������������������������������������������������� �����?������������        � �� � ?��� ��        p ����������?�>�y���}��������??�������������������������������������������������������������?�>�y���}��������??������������       ��ǁ�� ����?��        p ����������?�8~9���<��~���>�������������������������������������������������������������?�8~9���<��~���>������������       ����~ ������a�        p ������������ �?���9��>������������������������������������������������������������������ �?���9��>���������������        �o���=� 8�7c��         p �������������D�~��q��|��<Ȝ|<�����������������������������������������������������������������D�~��q��|��<Ȝ|<�������������        �o��8q� 1�>��         p �������������	��s��sǎ|��|�<�|�����������������������������������������������������������������	��s��sǎ|��|�<�|�������������        �8�0� 3�|Ä         p �����������������������|�<{����������������������������������������������������������������������������|�<{��������������        3�q�80c<1�cy��         p �������������3�#��Ϝ��8����~������������������������������������������������������������������3�#��Ϝ��8����~��������������       �7�a�81�xc�<c�>         p �����������g�s������x�Ü������������������������������������������������������������������g�s������x�Ü����������������       0w�8pg�xg����         p �����������ψ�GǏ�y����9�|8����������������������������������������������������������������ψ�GǏ�y����9�|8��������������       0fð0�n������          p �����������ϙ�<O�����?9�<�<����������������������������������������������������������������ϙ�<O�����?9�<�<��������������       0�9�pa�|��<���          p ������������1�8����O3��~y�8�������������������������������������������������������������������1�8����O3��~y�8����������������       3�1�`g`�0���y�8         p ������������3�p�����3��y�y�������������������������������������������������������������������3�p�����3��y�y����������������       �?�0��~`�a���0<         p �����������c� ���p3���y������������������������������������������������������������������c� ���p3���y����������������       �`�@<�@a����         p �������������	��?���xg���>��������������������������������������������������������������������	��?���xg���>����������������                         �          p �����������������������������?����������������������������������������������������������������������������������?��������������                                    p �������������������������������������������������������������������������������������������������������������������������������                                    p �������������������������������������������������������������������������������������������������������������������������������                                    p �������������������������������������������������������������������������������������������������������������������������������           8                         p �������������������������������������������������������������������������������������������������������������������������������           p                         p �������������������������������������������������������������������������������������������������������������������������������           �                         p �����������������������������������������������������������������������������������������������������������������������������           �                         p ��������������?����������������������������������������������������������������������������������?�����������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������   ��              �   0     �   p �����������������������?���������� ���������������������������������������������������������������������?���������� �������  �� �            �8   0    �   p �����>?�����������������?���������� ���������������������������������������������������>?�����������������?���������� �������  ��           0  �0   `        p �����|��������������������������������������������������������������������������������|������������������������������������                �0   �        p ���������������������������������������������������������������������������������������������������������������������������             8    |`   �        p ������������������������������ ���������������������������������������������������������������������������������� �������������  >            0    ?�`  �    �   p ����������������������������� �������������������������������������������������������������������������������� ������������  �< ��!� ��� � ? � �p ?�   p �������?�?�q����~�=����=���?����������������������������������������������������������?�?�q����~�=����=���?������������  �~1�`w���� �<  �  ?� 88   p �������?��?� ����|�<����0��������������������������������������������������������������?��?� ����|�<����0����������������  ��1�`�����`�x �3  s�     p �����O��?���b�q��y����a������g������������������������������������������������������O��?���b�q��y����a������g����������  >1�c�a���0s11���� �c  �     p ������9��'?�ό��c�x'���I�������������������������������������������������������������9��'?�ό��c�x'���I����������������  a�g c���0�cs0�� l�  �8     p �����y���F�8����?��O�������<��������������������������������������������������������y���F�8����?��O�������<������������   �� c7 �a��nq�0 0C�� �0     p �����<�8�����y�y?��?����ϼ3#���|��������������������������������������������������������<�8�����y�y?��?����ϼ3#���|������������   �� f~ g���` 0�� 9�8`     p �����<�1�������?����f���yǟ������������������������������������������������������<�1�������?����f���yǟ����������  �� lx f��À` 3�� �0�     p �����y�a�������<����x�����?������������������������������������������������������y�a�������<����x�����?����������  �� |� 8�?�� � g; �q�     p �����y�A��=���3��zx����������<�?������������������������������������������������������y�A��=���3��zx����������<�?����������  ;| x� ��{	�� 8� |3 g   0   p ������ă��9��'��pp���?�����������������������������������������������������������������ă��9��'��pp���?��������������������  s� p� ���� 0� �38 >8�   p   p �������3��1��?&$�`����?�����������������������������������������������������������������3��1��?&$�`����?�������������������  � `� �����> a� �c� 8�� �   p ������g����~`d���������������������������������������������������������������g����~`d������������������  � `p �1��� !� @a� �� �   p ������=�������p��������?����������������������������������������������������������=�������p��������?�������������          8                  � �    p ��������������������������������?�� �������������������������������������������������������������������������������?�� ��������          0                  �  �    p ���������������������������������������������������������������������������������������������������������������������������          p                  �       p �����������������������������������������������������������������������������������������������������������������������������          `                          p �������������������������������������������������������������������������������������������������������������������������������          �                          p �����������������������������������������������������������������������������������������������������������������������������          �                          p ������������?����������������������������������������������������������������������������������?�������������������������������         �                          p ������������?����������������������������������������������������������������������������������?�������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������   ��                     0           p ����������������������������������������������?�������������������������������������������������������������������������������   ��     �         0     0           p ����������������������������������������������9?�����?�������������������������������������������������������������������������   ��     �         0     0           p ����������������������������������������������9?�����?�������������������������������������������������������������������������   ��8�|��f�����9�sǏ9�6y��Ǐ9�   p ����������������������������������������������90���c�a���8p�Ɇd~8p��������������������������������������������������   �كm�3v���f��m�30flٳ06͛lٳ0   p ����������������������������������������������&|�g̉3'�L�?�g�ϙ�&L��2d��&L��������������������������������������������������   �ߟ1�?f���f���m�30g��06͛���   p ����������������������������������������������? `���0'�L�?3��Ϙ�L��2d�s�L�������������������������������������������������   ��3�0f��f�͛m�30f�06͛ ��    p ����������������������������������������������?'��ϙ3��L�?2d��ϙ��L��2d�3�L��������������������������������������������������   �ٳm�3f��3n�͛m�30flٳ0ͻlٳ0   p ����������������������������������������������?&L�g̙3'�̑?2d�g�ϙ�&L��2D��&L��������������������������������������������������   ��8�fg�>���l��cǏ1�x�Ǐ1�   p ����������������������������������������������?0��ᙘg���?3���8p���8p��������������������������������������������������                                    p �������������������������������������������������������������������������������������������������������������������������������                          p          p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������    ?�����������������������������    p �������                            �������������������������������������������������������������������������������������������    ?�����������������������������    p ������������������������������������������������������������������������������������������������������������������������������    ?�����������������������������    p ������������������������������������������������                           ��������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    8                           �    p ������������������������������������������������������������������������������������������������������������������������������    ?�����������������������������    p �������                           �������������������������������������������������������������������������������������������    ?�����������������������������    p ������������������������������������������������������������������������������������������������������������������������������    ?�����������������������������    p ������������������������������������������������                            ��������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������              �o߿   ` 6          p ������������������������������������������������������������� @���������������������������������������������������������������             c1�  ` 0 �        p ���������������������������������������������������������������|�������������������������������������������������������������             c1�  ` 0 �        p ���������������������������������������������������������������|�������������������������������������������������������������        3�9�c1���6��        p ������������������������������������������������������c��q����|a�p�������������������������������������������������������        6��6��c?3lٶ홀        p ������������������������������������������������������'�L�$�0�������&If������������������������������������������������������        3���1�3o�6���        p ��������������������������������������������������������L�����|���'�2������������������������������������������������������        �1����1�3l6́�        p ����������������������������������������������������$�g�L�y����|�����2~������������������������������������������������������        �v��6��1�3lٶ͙�        p ����������������������������������������������������$�'�L�$����|���&I2f������������������������������������������������������        q�1��c����6��        p ����������������������������������������������������s��q���N~a�p�3������������������������������������������������������                          �        p ������������������������������������������������������������������������������������������������������������������������������                                   p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p �������������������������������������������������������������������������������������������������������������������������������                                      p ���������������������������������������������������������������������������������������������������������������������������������������������������������������������� ��                                      ?����������������������������������������������������������������������������������������������������������������������������� ����������������������������������������������������������������������������������������������������������������������������������������������������������������������� �������������������������������������������                                       ��������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         �������������������������������������������������������������������������������������������������������������������������������                                         ������������������������������������������������������������������������������������������������������������������������������