�i  X  ��������������������������p��p��p��p��0��0��0��0������������������0��0��0��0� p� p� p� p� �� �� �� ������������������������������������������?��?��?��?��������������������������������������������������������������������� �     �    �    <    �    �    �                            �   � � � @ � � @ � �   .� 1� ?� @ ]  c� @ � �  ǀ �� 9 t � �  r �  �  � � < � � � x � � @ � �   .� 1� ?� @ ]  c� @ � :  G� ~� 9  4    =  2                                           ��< '� �  >���   ��? � ? �� 