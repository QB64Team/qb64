��a  �5w                            0           �                                                         0           �                                                         0           �                                                         0           �                                                         1�       � �                                                         1�       � �                                                         1�       � �                                                         1�       � �                                                         00       � �                                                         00       � �                                                         00       � �                                                         00       � �                                                         0><x��x<y��6�                                                         0><x��x<y��6�                                                         0><x��x<y��6�                                                         0><x��x<y��6�                                                         0;fͶ`f��6ـ                                                        0;fͶ`f��6ـ                                                        0;fͶ`f��6ـ                                                        0;fͶ`f��6ـ                                                        03f���|~}��6߀                                                        03f���|~}��6߀                                                        03f���|~}��6߀                                                        03f���|~}��6߀                                                                                                                                                                                                      03f�f �`̀f6�                                                                                                                                                                                                                                                                              1�fͶ`�f́�ـ                                                                                                                                                                                                                                                                             3<x��|<|���6�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   p                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �                                                                                    <                                                                                                                                                                                                     �        p    8                                                                 p    G                                                        @        p                                                                      p                                                            �        p    ~                                                        �        p    ��                                                                `                                                                      `                                                            �        p    ��                                                      �      p    `                                                                `                                                           �        `                                                             ��      p    �                                                      p      tp   �                                                                `                                                                      `           ?�  �      �   �                             ?�      p    �                                                      �     �p    `                                                                `                                                                    `           � ��      �� ?��                             ��     �p    �                                                      8�    � p    �     ?�  �      �   �                                       `                                                                   `            ������      ������                             ���    ��p    ��                      @                              �  ��p     `     � ��      �� ?��                                       `                                                                    `           ������      �����p                             ���  ���p     �     d    H      @   �                              � ��@ zp    �    ������      	?����`                                       `                                                                  � `           ������      ������                              {�������~p     �    0C    0      0                                       �p     p   �������      ������                                       `          @                                                     @� `            �?���?      ����s�                              ������p     �   � �  �       �   �                               �    �p     �   �?���>      ����s�                                       `                         �                                        @  `            �����      �w���      �  �      �   ?�     �����~p     ��  � x�        G� q                               �  ��p      p  p?����      �p���                                       `                                                                     `            ���}W�      ��7��      ?� ��      �� ��     ���  ?~       ?�  o� |��        w�*��                               �����      ���oȃ|W�      ��7�@      �  �      �   ?�             �       @                                                                        �����      ���?��      �����      ������      w���߿�|       � ��  |         @�                                 @@�       ` �� �����      ���?��      ?� ��      �� ��             �                        @                                                  �   �����      ����P      �����ۀ     ������      ���߿���      �����            A �      2    $          @         @@            ����      ����@      I�����      ������            ��                       @                                                 �  ?����      ����P      �����     �����x      ���߿��        �����@           �      !�            �          @             ����      ����@      ^����      �����p           @C�                                                                             ����       ����@      �������     ������      �������        ~����@            (�       `  `       F   F                     � @ ����        ���@      ����      ������         @@A�                                                  @                               �����       ����@      �ÿ�|�     �;����       �����         ��� �          �((*�       <@ ��       #� 8�                      a� ����        ���       Å�|      �8_���         @@                                                         �                           ? ����      ����       �A����     ����       �����         ���               ,(
�       �AT        ;�HP                        ��      ���       7�A�+�      ~D⿠           @                                                                                   ? ���      �M��       ?��A���      �����       �����         ���     2         ,�+"�         �          �                         ���        M��       �WA��       ��t��                                                                                                 ��       � �0       ������      �����       �����          }��              ,�)�                     �P                      � 	            �           ����       7����                                                                                                � �        < ��       ������      �����        ���           ��               ,� 
�                     �P                       b @           $            �����       �{���                                                                                                   �            �        ������      �����                       ��     3�        �#8                        	P                         �          	   �        7����       ���                                           0                                                      <  #�       � 8        ?����       ���j�                       ��               ��                      �P                         $           @           ����        ���j�                                                                                                              � �        ����        >��*�                        ~�                �                       T �P                       �  	            �           ���        ��*                                                                                                    �          < �        ����        ��.                         �     3�          8                      VR�P                        `   @          $  �         g���        )�(                                            0                                                       � #�         8         ���        ��(                         �                �                      R�P                            �           	            ��          ٭                                                                                                      <          ��         ��          9��                         �                                        RUP                        @   $           @                                                                                                                                           ��                      �                                3�          8           �         S=P                        �   	           � �                       �                                            0                                                      �#�         <8           "�          (                                           �                      �@                             @           $                                                                                                                                 ���         ��            @                                                                   ��          �@                              �                                                                                                                                            ��         ��          ��          �                                                          @           @                              ��         ��                                                                                                                                +�          �           +�          �                                           p                      p                                            �                       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ?0           ��       ?0           ��       >            >`                                                                                                                                                                                                                           1�          3` ��       1�          3` ��       3            c`                                                                                                                                                                                                                           1�          0` ��       1�          0` ��       3            ``                                                                                                                                                                                                                           1���        0vgϞ>       1���        0vgϞ>       3<����       `|y���                                                                                                                                                                                                                       ?0m�        flٳf       ?0m�        flٳf       >��`       `v͛6l                                                                                                                                                                                                                       03�        flٿf       03�        flٿf       3>��3�       `f͛7�                                                                                                                                                                                                                       06m�        flٰf       06m�        flٰf       3f͛6`       `f͛6                                                                                                                                                                                                                       06m�        3f�ٳf       06m�        3f�ٳf       3f͛6`       cf͛6l                                                                                                                                                                                                                       03�        3�Ϟ>       03�        3�Ϟ>       >>��3�       >fy���                                                                                                                                                                                                                                                                                        �                                                                                                                                                                                                                                                                                          �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          �                                                                    �                                                                                                                                                                                                                  �                                                                    �                                                                                                                                                                                                                  �                                                                    �                                                                                                                                                                                                                  �                                                                    �                                                                        |���  `ll             |���  `l          � 0`   �                                                                                   �                                                                    �                                                                        ���0  `�`             ���0  `�          � 0`   �                                                                                   �                                                                    �                                                                        ���   `�`             ���   `�          � 0`   �                                                                                   �                                                                    �                                                                        �σϏ`�l��             �σϏ`�6�        ͙����ǜ�                                                                                   �                                                                    �                                                                        �ف�nٳ`�훳             �ف�nٳ`���        ��6f��`��                                                                                   ����            ���     ���            ?���                          ����            ���     ���            ?���                              �ـ6ٳ`�m�3             �ـ6ٳ`���        ͛6f�����                                                                                                                                                                                                                                     �ـ6ٳ`�m�3             �ـ6ٳ`���        ͛6f�f��                                                                                                                                                                                                                                     �ك6lٳ`�m�3             �ك6lٳ`���        ͻ6c��l��                                                                                                                                                                                                                                     |ρ���`�l�3             |ρ���`���        ���� ����                                                                                                                                                                                                                                             �                      �                 �                                                                                                                                                                                                                                             `�                     `                �                                                                                   