�i  8���                      x      �                                                x      �                                                x      �                                                x      �                                                � � 0  �  �                                             � � 0  �  �                                             � � 0  �  �                                             � � 0  �  �                                             � � 0  �  �                                             � � 0  �  �                                             � � 0  �  �                                             � � 0  �  �                                             ��<y��9���8���                                            ��<y��9���8���                                            ��<y��9���8���                                            ��<y��9���8���                                            y�f̀37lٰ6��0                                            y�f̀37lٰ6��0                                            y�f̀37lٰ6��0                                            y�f̀37lٰ6��0                                                                                                                                                                  �~���3�l߰���                                                                                                                                                                                                                             �`���3l�0��                                                                                                                                                                                                                              ͛f́�36lٰ6Û0                                                                                                                                                                                                                             x�<x��1�g�0c��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �             ?��  ?��                                                   �   �                                     �             <�  <�                                    ` 0           � 0  � 0                ?�                 ���           ��� ���                                    ��           ���  ���                ?�                 �                                � �                                             �  ���                ����          ?��� ����              ���                ���           ��� ���           �    0                   �                �          � �                    �@           �   @@   @         ��� ?���             �  � ��         ����������          ��� ���                ?����          ���������           8                 �  @�@              �                 �?� �            ��             � 
 �          ��������           ���?���         �� ���� ��         ��� �����            �������         ����������           � ?� @             0�             �  �           ?� �� �           �   `          � �� �        �������          �������          ������         ���������            �����          ����������        �?� (� �            �            � �� �         � �p             <  x�� �          <  ��  ��       ��������          < �����         ���������       ����������            ?�����           ?�����������       � �p              @x �            @<  �|  �@        `  �   ��         �   � `         ��   `    `        ?���������         � ?����� `        �?����������       �����������           �����           ������������       0`  �   �                          �   `   `       C    � ?�             d��          �  �         �����������          �����         ������������       ����������           �����          ������������       �    ��                b                             ?� G���          ���         ������      ������������          �����         ������������       ������������           ����          ������������                          � @                         0�������        `  �_�   �        ��� ���� �      �����������|        `  �����  �       ����������      ������������           ����           ������������       0       �              �                 �    �      �?��������b        �  ����            ������`����`      ?����������        �  ���           ??������������     ������������           ����           ?������������       �    �    `            �            �     `    `�     �����a����           �k�          A��������@     ������������          ����          ��������������     ������������            ���           �������������           b    �           � d            �                ��������           ���          ��������      ������������          ����         ��������������     ������������           ����           ��������������        x      @           0                           �  ����          �	�          ?����������      �� ���������         ����         ��������������     �� ���������          ����          ��������������        0                                             � � ���      0     ǀ   �      ����������       �� ��������      0   ����   �     ��������������      � ��������          ���          ��������������      �`   8              �@                         @   ��  ��P      @    ���     @       �������������     @?  ���� ���      @   ���    @     ������������|        ���� ���          ����          ��������������      #       `  @          �                   �    �     �    ��� ��       �    ���           C�������@����@     �   ���p ���      �   ���p          ��������������         ���� ���          ����          ��������������             �                �          @       A    @         ��@  �         ��@          �������� ���         ?���� ���         ����         ?�������������         ?����  ��          ����          �������������             @ �               H           �        �            @?��   �	         $�~          !������������       ����  ?��         ;����         >��������������        ����  ��          ?���          ?���������������                            �$                  @            ��  ��        @?�?         @������A���@       �����  ���        ��?�         ��������������        ����  ���         ��?�          ����1����������        �                                 N               ��?	  ��@        ���         �?��  ��� ���        ���?�  ���        ����         �����������?����        ���?�  ���         ����          ���� ���������                             	              ��`              ����  ��          ���          ��  s��� ���       ����� ���       �����        ��������������       �����  ���         ����          ���� ����������          @                �                         � �@  �        ���        ���� ���� ���      �� ��  ��       �����        ��������������       �� ��  ��        �����         ���������� ����                                                         � �   ?�        � �@    �    A��� ���� ?��       �� ��  ?�p        �� ��    �    ��������� ���       �� ��  ?��        �� ��         ��������� ?���                �                         @  @   @     @    � �   �@    @    �  �     @    !��  ����� ���   @   �� ��  ��    @   �� ��    @    ?�� �����| ��|       �� ��  ��        ��  ��         ?�� ������ ���               @                               �    �   @    � ��  �    @   �  x�    @    S�� ����D ��D   @   �� �p  ��    @   ��  �p    @    _�� ������ ���       �� ��  ��        ��  �         �� ������ ���            �                  ��                 @   @   �   �  �H  �     �    �  |P         ���  ����@ ��@   �   ��  ��  ��    �   ��  �         ��� ������ ���       ��  ��  ��        ��  �         �� ������ ���            @                 @                 B    B       ?�  |    ~�        �  >         � ����" ��"      ��  �   ��       ��  ?�       �� ������ ���       ��  �   �        ��  ?�          � ������ ���                 �                         �0    
               �  <             �  (            ����  ��      ?��  ?�   >       ��  �        ?� ������  ���       ?��  ?�             ��  �             ������  ���             $   >                         ?�                �  >            ?�             ���  �      ��  ?�           ��  �           ������  ��       ?��  ?�             ��  �             �����  ��       @                                        �            �               ?�  �            ��?�  ?�      ��  �           ?��  �           ?������ ?���      �   �             ��  �             ���?��  ?��         �                                      @@ �   �      �               �  �            ?� ��� ���     ��   �           ?��  �           ?���?��� ?���      �   �             ?��  �             ?�� ��� ���      �                        
                �            �   �               �            ?� ��  ��      ��   �           ?�   �           ?�� ��� ���      ��   �             ?�   �             ?�� ��� ���            	                                               �   �           @�   �            � ��  ��     ��   �           �   �           �� ��� ���      ��   �             �   �             ?�� ��� ���                                           @    @   @    �   �            �   �           @� ��@ ��@    ��   ��          �   �           �� ��� ���     ��   �             �   �             �� ��� ���            �                                           �   �           �   �            � ��  ��     ��   ��          �   �           �� ��� ���     ��   ��            �   �             �� ��� ���                                                         �   �           ��   �            �� ��  ��     ��   ��          ��   ��          ��� ��� ���     ��   ��            ��   �             �� ��� ���                              �            �             �   �@          �    �          ��� ��  ��     ��   ��          ��   ��          ��� ��� ���     ��   ��            ��    ��            ��� ��� ���                                                        �   �           �    �            �  ��  ��     ��   ��          ��    ��          ��  ��� ���     ��   ��            ��    ��            ��  ��� ���                                                        �    �           �    y           �  ��  ��     ��   ��          ��    ��          ��  ��� ���     ��    ��            ��    �            ��  ��� ���                             �@                          �    �     �             y@    �          �� ��     ��   ��    �             ~�    �      ��  ��� ���     ��    ��                  �            �   ��� ���                                          �               �    ��    �             x�    �           ��  ��     ��    �`    �             @    �      �   ��� ���     ��    ��                  �           �    ���  ���            �                   �                           �    x�    �             <�    �          ��   ��      ��    �`    �             @    �      �    ���  ���     ��    �                  ?�           �    ���  ���            ��                  @�                             �    x�    �             <�    �            �   �      ��    �p    �             `    �      �    ���  ���     ��    �                  ?�           �    ��  ��            ��                  @�                �  �            x�    �             <�    �           �  �            p    �             ?`    �      �    ���  ���            �                  ?�           �    ��  ��             �                   �                 �   �  @          x�    @  @    @     <�    @  @         ��  �� @          p    @  @    @     ?`    @  @   �    �x  ��x            �                  ?�           �    ��  ��             �                   �                  �  � � @          x�    @  @    @     <�    @  @        ��  �� @          p    @  @    @     ?`    @  @   �    �|  �|            �                  ?�           �    ��  ��             �                   �                   �    � @    @     <@    @  @    @     @    @  @        ?��  ?�� @    @     �    @  @    @     ?�    @  @   �    �|  �|            ?�                  �           �    ?��  ?��            @@                   @                 @ �  @ � @    @     <@    @  @    @     @    @  @         ?�B  ?�@ @    @     �    @  @    @     ?�    @  @   �    ?��  ?��            ?�                  �           �    ?��  ?��            @@                   @                  @    B @    @     <@    @  @    @     @    @  @         �!  �  @    @     �    @  @    @     �    @  @   �    ?��  ?��            ?�                  �           �    ��  ��            @H                   @                       ! @    @     <@    @  @    @     @    @  @         �� � @    @     ?�    @  @    @     �    @  @   �    �� ��           ?�                  �           �    ��� ��             H                   @                     �@    @     <H    @  @    @     @    @  @         �� � @    @     ?�    @  @    @     �    @  @   �    ��� ���           ?�                  �           �    ��� ���            @                   @                      @    @     <H    @  @    @     @    @  @         ��  �� @    @     ?�    @  @    @     �    @  @   �    ��� ���           ?�                  �           �    ��� ���            @                   @                        @    @     <@    @  @    @     @    @  @          ��   �� @    @     ?�    @  @    @     �    @  @   �    ��� ���           ?�                  �           �     ��   ��             @                   @                  �  �@    @           @  @    @           @  @                  @    @           @  @    @           @  @                                                                                                                                        @    @           @  @    @           @  @           @      @    @           @  @    @           @  @           @                                                                                                                            @    @           @  @    @           @  @    @      @    @ @    @           @  @    @           @  @    @      @    @                                                                                                                       @    @      @    @  @    @      @    @  @    @      @    @ @    @      @    @  @    @      @    @  @    @      @    @                                                                                                                                   �    �              �    �              �    �             �    �              �    �              �    �                                                                                                                                   �    �              �    �              �    �             �    �              �    �              �    �                                                                                                                                   �    �              �    �              �    �             �    �              �    �              �    �                                                                                                                                   �    �              �    �              �    �             �    �              �    �              �    �                                                                                                                                   �    �              �    �              �    �             �    �              �    �              �    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �    �              �    �              �    �             �    �              �    �              �    �                                                                                                                                   @    @    @    @    @    @    @    @    @    @    @    @   @    @    @    @    @    @    @    @    @    @    @    @                                                                                                                         @    @    @    @    @    @    @    @    @    @    @    @   @    @    @    @    @    @    @    @    @    @    @    @                                                                                                                                   �    �              �    �              �    �             �    �              �    �              �    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �    �              �    �              �    �             �    �              �    �              �    �                                                                                                                                   @    @  @    @      @    @  @    @      @    @  @    @     @    @  @    @      @    @  @    @      @    @  @    @                                                                                                                           0    0 �   �      0    0 �   �      0    0 �   �     0    0 �   �      0    0 �   �      0    0 �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �    �              �    �              �    �             �    �              �    �              �    �                                                                                                                                   `    `�    �        `    `�    �        `    `�    �       `    `�    �        `    `�    �        `    `�    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �   `�   `          �   `�   `          �   `�   `         �   `�   `          �   `�   `          �   `�   `                                                                                                                               <  �<  �          <  �<  �          <  �<  �         <  �<  �          <  �<  �          <  �<  �                                                                                                                               � � � �           � � � �           � � � �          � � � �           � � � �           � � � �                                                                                                                                 �   �             �   �             �   �            �   �             �   �             �   �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     � �              0    `               �6                                                                                                                                                                                                6 �              1�    `                6                                                                                                                                                                                                 �              00    `                6                                                                                                                                                                                                <y�              0><����               �                                                                                                                                                                                                �f��              0;f͛6`               ��                                                                                                                                                                                                 6f��              03f͛�`               �                                                                                                                                                                                                 6f��              03f͛`               �                                                                                                                                                                                                6fͰ              1�f͛6`               �                                                                                                                                                                                                �<y�              3<����               �                                                                                                                                                                                                                      ��                                                                                                                                                                                                                                          ��                                                                                        