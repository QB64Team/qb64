�f  0�;L                                                       ��������������������                   ��������������������                                                           ��������������������                                                                                               ��������������������                   ��������������������                                                                                               ��������������������                   ��������������������                                                                                               ��������������������                                                         !���������������������                  !���������������������                                                        =                   �                  B��������������������@                  B��������������������@                  =                   �                  {                   �                  ���������������������                   ���������������������                   {                   �                  �                   �                 ��������������������                 ��������������������                  �                   �                 �                   �                 ��������������������                 ��������������������                 �                   �                 �                    �                 !��������������������                 !                   ?                 ����  ����   ����  �                 �                    |                 C���������������������                 B                   �                 ��m�$�H�m�ܒI$���m�$�|                 x                    >                 ����������������������                 �                   �                 {���  ����   ����  >                 �                                     !����������������������                !                   ��                ����  ����   ����                   =�                    �                B���������������������@                B                   �@                =�$�6�m�$�I#m��rI$�6�l�                {�                    �                �?���������������������                 �                    �                 {�  ���   ����   ���                ��                    �               ���������������������               @                    �                ��  ���   ����   ���               �                     �               ����������������������               �                    ~               �I$�6�m�$�I#m��rI$�6�m��               �                      �               !����������������������               !                     ?               �   ���   ����   ����               �                      |               C�����������������������               B                     �               �   ���   ����   ���|               x                      >               ������������������������               �                     �               zI$�6�m�$�I#m��rI$�6�m�>               �                                     !������������������������              !                     ��              �   ���   ����   ���               =�                      �              B�����������������������@              B                     �@              =�   ���   ����   ����              {�                      �              �?�����������������������               �                      �               {�I$�6�m�$�I#m��rI$�6�m��              ��                      �             �����������������������             @                      �              ��   ���   ����   ����             �                       �             ������������������������             �                      ~             �`   ���   ����   ����             �                        �             !������������������������             !                       ?             �rI$�6�m�$�I#m��rI$�6�m� �             �                        |             C�������������������������             B                       �             ��   ���   ����   ��� |             x                        >             ��������������������������             �                       �             {�   ���   ����   ��� >             �                                     !��������������������������            !                       ��            �rI$�6�m�$�I#m��rI$�6�m�              =�                        �            B�������������������������@            B                       �@            =��   ���   ����   ��� �            {�                        �            �?�������������������������             �                        �             {��   ���   ����   ��� �            ��                        �           �������������������������            @                        �             ��rI$�6�m�$�I#m��rI$�6�m�$�           �                         �           ��������������������������            �                        ~            ��   ���   ����   ��� �           �                         �           !��������������������������            !                         >            ���   ���   ����   ��� �           �                         �           C��������������������������            B                                     ��rI$�6�m�$�I#m��rI$�6�m�$��           x                         �           ���������������������������            �                                     {��   ���   ����   ��� �           �                         �           !��������������������������            !                                     ���   ���   ����   ��� �           =�                         �           B��������������������������            B                                     =��rI$�6�m�$�I#m��rI$�6�m�$��           {�                         �           �?��������������������������            �                                      {���   ���   ����   ��� �           ��                         �          ��������������������������           @                                     ����   ���   ����   ��� �          �                          �          ���������������������������           �                                    �6�rI$�6�m�$�I#m��rI$�6�m�$��          �                          �          !���������������������������           !                                     ����   ���   ����   ��� �          �                          �          C���������������������������           B                                     ����   ���   ����   ��� �          x                          �          ����������������������������           �                                     zI$���m�$�H�m�ܒI$���m�$�H�m�          �                          �          !���������������������������           !                                     �  ����  ����   ����  ���          =�                          �          B���������������������������           B                                     =�  ����  ����   ����  ���          {�                          �          �?���������������������������           �                                      {�I$���m�$�H�m�ܒI$���m�$�H�m�          ��                          �         ���������������������������          @                                     ��  ����  ����   ����  ���         �                           �         ����������������������������          �                                    �   ����  ����   ����  ���         �                           �         !����������������������������          !                                     ޒI$���m�$�H�m�ܒI$���m�$�H�m�         �                           �         C����������������������������          B                                     �   ����  ����   ����  ���         x                       �  �         ����������������������������          �                       �            x   ����  ����   ��������         p                       �  �         �����������������������������          �                       �            t�I$���m�$�H�m�ܒI$���m�/�H�m�         `                       �  �         ����������������������������          �                       �            h   ����  ����   ��������         @                       �  �         ����������������������������          �                       �            X   ����  ����   ��������                                 
  �         ����������������������������          �                       ;�            �I$���m�$�H�m�ܒI$���m�?�H�m�                                 ;�  �         �����������������������������          �                       4            x   ����  ����   ����?����                                 >>  �         �����������������������������          �                       0            x   ����  ����   ����>>���                                 <
  �         ����������������������������          �                       0            \�I$���m�$�H�m�ܒI$���m�<H�m�                                 8  �         ����������������������������          �                       0            x   ����  ����   ����8���                                   �         ����������������������������          �                                   x   ����  ����   �������                                 8  �         �������������������������#���          �                                   \�I$���m�$�H�m�ܒI$���m�>>H�m�                                 �  �         ����������������������������          �                       �            x   ����  ����   ��������                                 �  �         ����������������������������          �                       �            x   ����  ����   ��������                                     �         �����������������������������          �                                     \�I$���m�$�H�m�ܒI$���m�$�H�m�                                     �         �����������������������������          �                                     x   ����  ����   ����  ���                                     �         �����������������������������          �                                     x   ����  ����   ����  ���                                     �         �����������������������������          �                                     \�I$���m�$�H�m�ܒI$���m�$�H�m�                                     �         �����������������������������          �                                     x   ����  ����   ����  ���                                     �         �����������������������������          �                                     x   ����  ����   ����  ���                                     �         �����������������������������          �                                     \�I$���m�$�H�m�ܒI$���m�$�H�m�                                     �         �����������������������������          �                                     x   ����  ����   ����  ���                                     �         �����������������������������          �                                     x   ����  ����   ����  ���                                     �         �����������������������������          �                                     #m��rI$�6�m�$�I#m��rI$�6�m�$��                                     �         �����������������������������          �                                     ����   ���   ����   ��� �                                     �         �����������������������������          �                                     ����   ���   ����   ��� �                                     �         �����������������������������          �                                     #m��rI$�6�m�$�I#m��rI$�6�m�$��              p  �                 �         �����������������������������          �    p  �                           ���� p ���   ����   ��� �                                   �         �����������������������������          � >   �  �                           ���� � ���   ����   ��� �                                  �         �����������������������������          �   �  �                           #m��rI��6���$�I#m��rI$�6�m�$��                                  �         �����������������������������          �   �  �                           ����� ���   ����   ��� �                                     �         �����������������������������`         �   �  �                 `         ����� ���   ����   ��� �           @                       @         �����������������������������         �   �  �                  �         #m��rI��6���$�I#m��rI$�6�m�$�@           `  �                    >�         �����������������������������          � _  |  �                 A          ����� ���   ����   ��� >�           `  �                    }�         ����������/������������������          � _  |  �                 �          ����� ���   ����   ��� }�           `  �                    ��         ����������/�����������������          � _  |  �                          #m��rI��6���$�I#m��rI$�6�m�$��           `  �                   ��         ����������/�����������������          � _  |  �                          ����� ���   ����   �����           `  �                   ��         ����������/�����������������          � _  |  �                          ����� ���   ����   �����               �                   ��         ����������/�����������������           � _  |  �                           #m��rI��6���$�I#m��rI$�6�m�'��               �                   ��         ����������/�����������������@          � _  |  �                @          ����� ���   ����   �����               �                   �         ����������?������������������          �    x  �                 �          ���� � ���   ����   ����                                    >��         ����������?�����������������           �    p  �                A           #m��rIt�6��$�I#m��rI$�6�m�>��                                    }��         ����������������������������           �                          �           ����   ���   ����   ���}��                                    ���         ���������������������������           �                                    ����   ���   ����   ������                                   ���         ���������������������������           �                                    #m��rI$�6�m�$�I#m��rI$�6�m����                                   ���         ���������������������������           �                                    ����   ���   ����   ������                                   ���         ���������������������������            �                                     ����   ���   ����   ������                                   ���         ���������������������������@           �                         @           #m��rI$�6�m�$�I#m��rI$�6�m����                                   ��         ����������������������������           �                          �           ����   ���   ����   �����                                   >���         ���������������������������            �                         A            ����   ���   ����   ������                                   }���         ���������������������������            �                         �            #m��rI$�6�m�$�I#m��rI$�6�m}���                                   ����         ��������������������������  @         �                          @         ����   ���   ����   ������                                  ���          ��������������������������  �         �                          �         ����   ���   ����   �����                                   ���          ��������������������������           �                                   \�I$���m�$�H�m�ܒI$���m�$����                                   ���          ��������������������������            �                                    x   ����  ����   ���� ���                                   ���          ��������������������������@           �                        @           x   ����  ����   ���� ���                                   ��          ���������������������������           �           ��������������           \�I$���m�$�H�            ��                      ����������������          �������������                        �                                   x   ����  �����������������                      ����������������          �������������                         �                                    x   ����  �����������������                      ����������������          �������������              @          �                         @          \�I$���m�$�H�����������������                                  ��           ��������������������������  �          �           �������������  �          x   ����  �            ��                                   ��           ��������������������������            �           �������������            x   ����  �            ��                                   ��           ��������������������������            �           �������������            \�I$���m�$�H�            ��                   ��             ��           ���       ?���������������            � �������� �������������            x ���������            ��                   ����            ��           �           �������������            ��������������������������            ������������            ��              �����������           ��                    ������������            ���������������������������            ����       ?���           ��            ?��������������          ��               0     �����������            ����������������������������            ���           ��          ��           �����������������         ��              @`     ���������� @         ?���������������������������� @         ?�              ��         ��          ������������������         �              @  @     ���������� �        �����߿�߿������������������� �        �                �         �          ?�������������������        �          
0 @     �  � ?���������         ���������������������������         �                 �        �         ��������������������        �                 �P       ���������         ?��������O��������������������         <                  �        �         ��������������������        �             @ � 	  @   ���������         ?����������������������������                                      �         ?��������������������        �            @H        
  0���������         ?�����������������������������                                      �         ?��������������������        �                � @ B ����������         �������������~���������������         �                           �         ?��������������������        �          @@ B      !  ��������         ?������������������������������         ?�                   �       �         ���������������������       �            &   @� �    � ��������@       �����������?�������z����������@       �                    �       �        ?�����������������������                  R     D   @     ���������       �������������������������������       ��                     �              ������������������������               �    �   � �������       ��W���������������{������������       �                       �              �������������������������                 �      $@   ��������       ����������������ۿ������������                                            �������������������������                � 	     �@ @�P   H �������       ��_������������/���������������                                               �������������������������                    �          � �������       �������������������~�����������                                               �������������������������               �   @� � �    �  D              }������n���7������������                                     �             �������������������������               � @  @     @  @                  ��߿����������������������            �                        �             ��������������������������                   �
@  �� J  
  @�               ?�������O������������?����           ?�                         ?�           ���������������������������              @  @P    ��  `                 ����߿���������������������          �                          �           ?����������������������������            4 %P  � � ��@                 ����������o������}�����������         �             �           �         ������������������������������                @   ��  ��   @              ������������������������������         ~          ��  ��          �         ������������������������������            �     @��� '���      @P         ������������������������������        �         ���  ���          |         ������������������������������          �    
  ����� ����    $           ������������������������������        �        ����� ����                 ��������������������������������                ������H������  0           ��������������������������������                ������ ������        �       ����������   ����  �����������        `  �  @�   ����  ��               ?���������   ����  �����������       8        �   ����  ��        �       ����������   ����   ����������        � ! �   ����   �  ! �         {���������   ����   ���������       `        �   ����   �        0       ?����������   ���    ����������        r @ ��   ���    �    P�@       �����������   ���    ���������       �       ��   ���    �               ����������   ���    ����������         H P@ �������������            �����������������������������       �       ������������               ����� ����  ���  � ���� ?����        � �����������������         ��������������������}�������           �� ������������� ��           ����   ����  ���  � ���  ����       @ ���@?�����������������@         ������������������������������          ��� ?����������������           ����   ���  ��� � ���   ���       ?����������������������� B        ��������������������?�����������          ?���������������?�������          ���    ���  ��� � ��    ���          �������������������������         ��������������������?�����������          ����������������?��������          ���    ��� > ��� � ��    ���       �� ?���������������������          ����� ?�����������������������         �� ?��������������������          ��    ���  p�� p  ?�� � ���         ��������������?�?��� ?��         ����������������?�?���������         ��������������?�?������          ?��  � ���   � �    ?�� �   ���         /��� ���� �� �� �?������          ?���������� ����� �?����������         �������� �� �� �?�������          ��   p ��� �� ?�?� �� p   ���        ����?������ ?�?���������         ������?�������?�?����������         ����?������ ?�?��������          ��     ������� ��� ���     ��        ������������� ���|������         ��������������������|���?�����          ������������� ���|���?���          ��     ��������������    ��         �����������������y�������C         �������������������y���������          ����������������y�������           �     ������� �������    ��          ������������ ��������������          �����������������?����������          ������������ ���?���������           �     ����� �������    ��           ������������ ���������?���           �����������������?�����?�����           ������������ ���?�����?���           ��   ����� ��������    �            ?����������� �������������           ����������������������������            ?����������� ������������            ?�   ������� ��������   ��            ����������� ������������             ?���������������������������            ������ ���� ����������             �   ������� ���������  �            ���������� ��������g���             ~��o����������������������              ���� ?��� ����� �����                  ������� ��������   �                  ������� ��������                     �����������������   �                  �� ��� ����� �                       ������  �������                       ������  �������                       ����������������                       � ?���  ������                       ?��� ?�� ������                       ?������� �������                       ?����������������                       ?� ����  ������                       ������ �� ����                       ������� �������                       ����������������                       ������  �������                       ������ �����                        ����� �   ����                        ���������������                        ������  ������                        ���?��� �����                        ������� ������                        ���������������                        ������  ������                         �����` ������                         �����` ������                         ��������������                         �����  ������                         �����P ������                         �����P ������                         ��������������                         �����  ������                         ����0 �����                          �����0 ������                         �������������                         ����  �����                          ���� �����                          ����� ������                         �������������                         ����  �����                          ����������                          ������������                         ��������������                         ����� �����                          �����������                          �������������                         ��������������                         ����� �����                             ���?��                            �������?������                         �  ���?��  �                         x  �� ?�� �                             �� ���                            ������ �������                         �  ������  �                         \�I?�� ���H�                             �����                            �������������                         �  �����  �                         x  ����� �                             ������                            ��������������                         �  ������  �                         x  ������ �                                                                ����     ?����                         �  ������  �                         \�I      $�H�                                                                ����     ?����                         �  ������  �                         x          �                                                                ����     ?����                         �       �  �                         x          �                                                                ����     ?����                         �       �  �                         \�I      $�H�                                                                ����     ?����                         �       �  �                         x          �                                                                ���������?����                         �       �  �                         x   ����  �                                                                ���������?����                         �       �  �                         \�I$���m�$�H�                                                                ��������������                         �           �                         x   ����  �                                                                ��������������                         �           �                         x   ����  �                                                                ��������������                         �           �                         \�I$���m�$�H�                                                                ��������������                         �           �                         x   ����  �                                                                ��������������                         �           �                         x   ����  �                                                                ��������������                         �           �                         \�I$���m�$�H�                                                                ��������������                         �           �                         x   ����  �                                                                ��������������                         �           �                         x   ����  �                                                                ��������������                         �           �                         \�I$���m�$�H�                                                                ��������������                         �           �                         x   ����  �                                                �              ��������������                         �           �         �              x   ����  �                                                �              ��������������                         �           �         �              #m��rI$�6�m�'                                                �              ��������������        �              �           �         �              ����   ���         �                                    �              ��������������       D              �           �         p              ����   ���        �                                 |  �              ��������������         �              �           �      |  �              #m��rI$�6�m�'          �                                 �  �              ��������������       0               �           �      �  �              ����   ���        0                                 �  �              ��������������       0               �           �     �  �              ����   ���        0                                 ��@�              ��������������       8b              �           �     ��@�              #m��rI$�6�m�'        8b                                ���                ��������������       8D              �           �     ���                ����   ���       (8D                                ��@               ��������������     @<H              �           �     ǀ@               ����   ���      x<H                                ��ǯ ?�            ��������������       <8P�             �           �     ǃǯ ?�            #m��rI$�6�m�'       8?���                               ��Ϯ �            ��������������       <0Q��             �           �     ��Ϯ �            ����   ���        ����                               �C V ��            ��������������      �0i�             �           �     �C  ��            ����   ���       �0?�                                �� � ��            ��������������      ~0��             �           �      ��   ��            #m��rI$�6�m�'      �0	�                                |  @ ��            ��������������     �~pH�	             �           �      |    ��            ����   ���      �~p�                                 �  ��            ��������������     O�|p��             �           �       �  ��            ����   ���      O�|p��                                � ��            ��������������     o�8<�            �           �       �  ��            #m��rI$�6�m�'      o�8<�q                                � �            ��������������     /�93���             �           �       �  �            ����   ���      /�83���                                 � ?�            ��������������    ��81Q�              �           �       � ?�            ����   ���     ��81Q�                                  � �            ��������������    ���q#              �           �       � �            #m��rI$�6�m�'     ���q3g �                             �    �            ��������������     ?���:~7             �           �    �     �            ����   ���      ?���:r7�                             � >   �            ��������������     ���<pn             �           �    �     �            ����   ���      ���<po�                             �     x            ��������������     ���4a�             �           �    `     x            #m��rI$�6�m�'      ����4a�x                             ��   <            ��������������     �����             �           �    �    <            ����   ���     >����<                             ��               ��������������     �����`             �           �    �                ����   ���     ����`                             �>   ?�            ��������������     ���#�J~            �           �     �    ?�            #m��rI$�6�m�'     ���#�J~                              �   ?�            ��������������    ����/�@            �           �           ;�            ����   ���     ���/�D                             �    ?�            ��������������     ǿ�?��`            �           �          ?�            ����   ���     ~��?��g                             8    p �           ��������������     ������            �           �    8      �           #m��rI$�6�m�'     8�������                            8    � �           ��������������     ?�������            �           �    8      �           ����   ���     8?�������                            p   p�  �           ��������������    ������            �           �    p   p   �           ����   ���     w����'.���                            p   ��  !�           ��������������    ��� ���            �           �    p   �   !�           \�I$���m�$�H�     w��� ���                            � �p  p�           ��������������    ��� |�             �           �    � �   p�           x   ����  �     ���� � �                            � �� � �           ��������������     ��S���             �           �    �  �    �           x   ����  �     �}�:S��x �                            � �� � �           ��������������     ��#����            �           �    � A�    �           \�I$���m�$�H�     ��:#��?��                           �@�� � �           ��������������     �����            �           �   �@ �   �           x   ����  �    �;����                              �p � p           ��������������   �������            �           �       p � p           x   ����  �    �;�����p                           � �  � p           ��������������   ������            �           �   � @    p           \�I$���m�$�H�    ��;���p                           � �  � 0           ��������������   ���������           �           �   �        0           x   ����  �    ���y���?��                           �    � 0           ��������������   ����� @           �           �   �       0           x   ����  �    	�����| p                           �    t|  8           ��������������   ����� H           �           �   �    |  0           \�I$���m�$�H�    ������ x                           �    .�  x           ��������������    ��� ��           �           �   �    �  p           x   ����  �    ���� ��x                           �p   �  x           ��������������    ��: �           �           �   �p   �  p           x   ����  �    ���: �x                           � � �� x           ��������������    ����            �           �   �    �� p           \�I$���m�$�H�    ���x�!x                           � � �� |           ��������������   �����D            �           �   �    �� p           x   ����  �    ���?��D |                           � � �� �           ��������������   ���� <            �           �   �    �� �           x   ����  �    �����8< �                           � ���� �           ��������������    ������            �           �    �   �� �           \�I$���m�$�H�    ����� �                           ����� �           ��������������    8��� �           �           �    �   �� �           x   ����  �    �8��8��                           ������ �           ��������������    p��XD?�           �           �    �� @�� �           x   ����  �    �p>NHD?��                           ����;���           ��������������   �r?��|@�           �           �    p� ����           \�I$���m�$�H�    �r<x�D@��                           �� �� �           ��������������   ����X �@           �           �    p� @� �           x   ����  �    ���XH �A�                           �    � �           ��������������   ���A �@           �           �    8    � �           x   ����  �    ���A �C�                           �     | �           ��������������   �w�A��            �           �    8     | �           \�I$���m�$�H�    ��A��#�                           �                  ��������������   � w��G��            �           �           �           x   ����  �    � w��G���                           �                  ��������������   � G��G�             �           �           �           x   ����  �    � G��G� �                           �                  ��������������   � ��@��            �           �           �           \�I$���m�$�H�    � ��@���                           �                  ��������������   � 9�P��            �           �           �           x   ����  �    � 9�P���                           ��     <           ��������������   � 8S��            �           �    �     ?�           x   ����  �    ��8S��?�                           �� �   x8           ��������������   �  0G�8 8           �           �    � �   �           \�I$���m�$�H�    �� 0W�8�                           �� �  �8           ��������������   �   o� 8           �           �     � �  ��           x   ����  �    ��  o�	��                           �� �  �8           ��������������   �  "n  8           �           �     � �  ��           x   ����  �    �� "n��                           �� �  �p           ��������������   ��   ,  p           �           �     | �  ��           #m��rI$�6�m�'    ��   ,��                           �� �  �p           ��������������   ��   (  p           �           �     > �  ��           ����   ���    ��   (��                           �π   > p           ��������������   �� 0 "  p           �           �     ?�   ?��           ����   ���    ���0 "?��                            ���    � �           ��������������    ��   $  �           �           �     �    ��            #m��rI$�6�m�'     ���  $���                            ���   ��           ��������������    ��   8 �           �           �     �   ��            ����   ���     ���  8���                            ���   ��           ��������������    ��   0  �           �           �     �   ��            ����   ���     ���  0���                            ��  � �           ��������������    �      �           �           �     ��  ���            #m��rI$�6�m�'     ���  ����              �����        ��  ��           ����    �����    �     �           �  �����   �     ��  ���            �����������     ���  ����                 �         ��� �x�           ����  � �����    ��    x�           �  ����   �      ?� ���            �����������     ��� ����                         ?��������           ����  �����    ?��   ��           �  �����   �     �����            #m��������m�'     ?���������                         ?�<����           ����  �����    ?�<   ��           �  �����   �     ������            �����������     ?���������                 �        ��  �             ����  ������    ��  �             �  ����   �      �����            �����������     ��������                  �        ��� � >            ����  ������    ��� � >            �  ����   �      |����            #m��������m�'     ��������                 p@        ����  ~            ���� p@�����    ����  ~            �  ��   �      ?�  ���            �����������     ��������                 �@        ����  �            ���� �@�����    ����  �            �  ����   �      � ��             �����������     ��������                 �@        ��    �            ���� �@�����    ��    �            �  ����   �      �����             #m��������m�'     ��������                 �@        ��    �            ����  �@�����    ��    �            �  ��G��   �      �����             �����������     ��������                 p@        ��    �            ����  p@�����    ��    �            �  �����   �      �����             �����������     ��������                  �         ���   ?�            ����   ������     ���   ?�            �  ����   �       ����             #m��������m�'      ��������                   �         ��   �            ����  ������     ��   �            �  ����   �       ?����             �����������      �������                            ?��  ��            ����  �����     ?��  ��            �  �����   �       ���              �����������      ?�������                            ��  �             ����   �����     ��  �             �  �����   �        ���              #m��������m�'      ������                   x          �����             ����  � �����     �����             �  �����   �        �               �����������      ������                              ������             ����    �����     ������             �  �����   �                         �����������      ������                               ������             ����    �����      ������             �          �                         #m��    �m�'       ������                                �����             ��������������      �����             �           �                         ����   ���       �����                                ����              ��������������      ����              �           �                         ����   ���       ����                                 ����              ��������������      ����              �           �                         #m��rI$�6�m�'       ����                                  ����              ��������������       ����              �           �                         ����   ���        ����                                  ��               ��������������       ��               �           �                         ����   ���        ��                                   ��               ��������������       ��               �           �                         \�I$���m�$�H�        ��                                                     ��������������                         �           �                         x   ����  �                                                                ��������������                         �           �                         x   ����  �                                                                ��������������                         �           �                         \�I$���m�$�H�                                                                ��������������                         �           �                         x   ����  �                                                                ��������������                         ��������������                                                               �������������                                       �                                      �                         �������������                          �������������                                       �                                      �                         �������������                          �������������                                       �                                      �                         �������������                                                                  ��������������                         ��������������                                                                                                         ��������������                         ��������������                                                                                                         ��������������                         ��������������                                                                                                         ��������������                         ��������������                                                                                                         ��������������                         ��������������                                                                                                         ��������������                         ��������������                                                                                                         ��������������                         ��������������                                                                                                         ��������������                         ��������������                                                                                                         ��������������                         ��������������                                                                                                         ��������������                         ��������������                                                                                                         ��������������                         ��������������                                                                                                         ��������������                         ��������������                                                                    ��������                            ���       ���                         ���       ���                            ��������                               ��������                            ���       ���                         ���       ���                            ��������                               ��������                            ���       ���                         ���       ���                            ��������                               ��������                            ���       ���                         ���       ���                            ��������                               ��������                            ���       ���                         ���       ���                            ��������                               ��������                            ���       ���                         ���       ���                            ��������                               ��������                            ���       ���                         ���       ���                            ��������                               ��������                            ���       ���                         ���       ���                            ��������                               ��������                               �                                      �                                      ��������                               ��������                               �                                      �                                      ��������                               ��������                               �                                      �                                      ��������                               ��������                               �                                      �                                      ��������                               ��������                               �                                      �                                      ��������                               ��������                               �                                      �                                      ��������                               ��������                               �                                      �                                      ��������                               ��������                               �                                      �                                      ��������                               ��������                               �                                      �                                      ��������                               ��������                               �                                      �                                      ��������                               ��������                               �                                      �                                      ��������                                                                       ���������                               ���������                                                                                                               ���������                               ���������                                                                                                               ���������                               ���������                                                                                                               ���������                               ���������                                                                                                               ���������                               ���������                                                                                                               ���������                               ���������                                                                                                               ���������                               ���������                                                                                                               ���������                               ���������                                                                                                               ���������                               ���������                                                              �     <  8   �                   sm�ܒI$���m�$p    � A������                  p            p    �  |   ��                  ��������������    � ��?���                  �            �       |   �                   w���   ���� p    � �������                  p            p    �� �   �                  ��������������    �  �|�@�                  �            �     � �   �                   w���   ���� p    �� �|�O��                  p            p    �� �   �                  ��������������    � �p� �                  ��������������     � �   �                   p            p    ���p���                  �������������    �� �   >�                  �                �  `� �                  �                 � �   ?�                   �������������    �� `�?��                  �������������    �� |   |�                  �                �  @� �                  �                 � |   �                   �������������    �� @���                  �������������    �| 8  ��                  �                � �� �                  �                 � 8  ��                   �������������    �������                                    �    �                   ��������������    �   �                    ��������������      �    ��                                     ��  ���                                     ���   �                   ��������������    ��  ��                    ��������������      �   ��                                     ��� ����                                     ���   ?                    ��������������    ��  �                     ��������������      �   ?��                                     ��� �?��                                     ��  �                    ��������������    ��                         ��������������      ?�  ���                                     ���  ���                                     ��  �p                   ��������������    ��     p                   ��������������      �  ���                                     ���  ���                                     ��� ���>                   ��������������    ��    �>                   ��������������      �� ��?�                                     ���� ����                                     ������<                   ��������������    ��   �<                   ��������������      �����                                     ���������                                     ������< |                   ��������������    ���   < |                   ��������������      ������                                     ���������                                      ��  � �                   ��������������     ��  � �                   ��������������      �����                                       ���������                                      �� ��                   ��������������     �� ��                   ��������������      ���?�                                       ��������                                      � ��� �                   ��������������     � ��� �                   ��������������      �  ��                                       ��������                                      ?� �� �                   ��������������     ?� �� �                   ��������������       �� ��                                       ?��������                                      ��    �                   ��������������     ��    �                   ��������������       �����                                       ��������                     ��������        ��    ?�                   ���        ���     ��    ?�                   ���        ���       �����                      ��������        ��������                     ��������        ��    �                   ���        ���     ��    �                   ���        ���       �����                      ��������        ��������                     ��������        ��   �                    ���        ���     ��   �                    ���        ���       ����                       ��������        �������                      ��������        ��   �                    ���        ���     ��   �                    ���        ���       ����                       ��������        �������                      ��������        ���  �                    ���        ���     ���  �                    ���        ���        ?���                       ��������        �������                      ��������         ��  ��                    ���        ���      ��  ��                    ���        ���        ��                        ��������         ������                      ��������         ?�����                    ���        ���      ?�����                    ���        ���         �                        ��������         ?������                      ��������         ������                    ���        ���      ������                    ���        ���                                   ��������         ������                      ��������         �����                               �        �����                               �                                     ��������         �����                       ��������         �����                               �        �����                               �                                     ��������         �����                       ��������          �����                               �         �����                               �                                     ��������          �����                       ��������          ?����                               �         ?����                               �                                     ��������          ?����                       ��������          ���                                �         ���                                �                                     ��������          ���                        ��������           ���                                �          ���                                �                                     ��������           ���                        ��������           ��                                �          ��                                �                                     ��������           ��                        ��������                                              �                                             �                                     ��������                                      ��������                                              �                                             �                                     ��������                                      ��������                                              �                                             �                                     ��������                                      ��������                                              �                                             �                                     ��������                                                                                     ���������                                     ���������                                                                                                                                   ���������                                     ���������                                                                                                                                   ���������                                     ���������                                                                                                                                   ���������                                     ���������                                                                                                                                   ���������                                     ���������                                                                                                                                   ���������                                     ���������                                                                                                                                   ���������                                     ���������                                                                                                                                   ���������                                     ���������                                                                                                                                   ���������                                     ���������                                      