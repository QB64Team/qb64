��^  H`�e                    �    �  m�`   ` �                                        �    �  m�`   ` �                                        �    �  m�`   ` �                                        �    �  m�`   ` �                                        0   �  l `� ` �                                        0   �  l `� ` �                                        0   �  l `� ` �                                        0   �  l `� ` �                                            �  l `� ` �                                            �  l `� ` �                                            �  l `� ` �                                            �  l `� ` �                                        ��������|�s�g�<y�p                                       ��������|�s�g�<y�p                                       ��������|�s�g�<y�p                                       ��������|�s�g�<y�p                                       �m�6 `�6m�v��l�fͳ`                                       �m�6 `�6m�v��l�fͳ`                                       �m�6 `�6m�v��l�fͳ`                                       �m�6 `�6m�v��l�fͳ`                                        7������m�f�co�`ͳ`                                        7������m�f�co�`ͳ`                                        7������m�f�co�`ͳ`                                        7������m�f�co�`ͳ`                                                                                                                                                                  6�`̓6m�f�3l`ͳ`                                                                                                                                                                                                                              6m�6`͛6m�f��l�fͳ`                                                                                                                                                                                                                              ���������f`q�g�<y�f�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          >   8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �        �                                                 |        �                                                 �        �                                                         �                                                 '�        #@                                                ?~        @                                                ?�        ��                                                                                                           �        ��                                                0_        ؠ                                                ?�        ��                                                `        ؀                                                ?�        �p          J�                                    ?'�       �p         ��                                    ?��       ��          ��                                    X        �`         B`                                    �@       !�         �       �           ��            w9�       �         ��       ��                         ��       ��         ��       �           ��       ��   HF        �          B       �           ��            ��        p         ��       ��          #         ���   w?�        p         E�       ��          <��       ���   ��       ��         ��       ��          ?��       �     H@         p         �       ��          !         �     x��       �         ��       �p          #         �    w?�       �         ��      �r          <��       ���   ��       ��         ���      ��          ?��       �     H@        �         G�@      �p          !         �     H��       ��         ��       ��          ?��       ���   w?�       ߘ         ���      ��                   ���   ��       ��         �?�      ��          ?��       ���   H@        ߘ         B       ��          =��       ���   _�p       p�         K�       	/v          ?��       ���   w��       p�         �<�      	v�                  ���   ~?�       ��         ���      ��          ?��       ���   H          �         @       	v          =��       ���   k��       �         O�      ��          #        �p   v?�       �         ��`      ؏�         <��       ���   }��       w�         ���      �          ?��       �     H                  A��      �          !         �     O�`       ��         O��      ��          #>        ��   u��       w�         �_`      �w          <��       ���   {��       ��         ���      ￀         ?��       �p    I�        s�         A@�      �7          !         �     O�        ��          O�      ��          #        ��   u_�       W�         ���      �          <��       �w�   {��       ��         ���      ￀         ?��       ��    I@        S�          A�       �?          !        �p    �`       ��          K�       ��                  ���   5��       w�         �/�      �q          ��       �W�   {��       ��         ���      ￀         ?��       ��    	�        s�          @#       �1                  �P    +��       �         ��       ��                  ���   6/�       �         ���      ؂          ��       �w�   }��       �         �{�      ���         #>       ��                       B       Ђ          ��       �p    �p       
v�          J,       /v          ;        ��   7��       
d�         ���      	F�         ��       ���   ~�       ��         J?�      ��          #       �|            
�         ��@      F          ��       �    ��       ��         J�       ��          �       �v   w�       Ґ         ��      �,          �~       ���   ?��       ��         J�       	?�          #�       �    H        Ҁ         ��      ,          �|       �    �        ��         �       �X          ��       ���   w%�       �l         ��       	            �       ���   �        ��         ��       ��          ?��       ���   8E�       �                  	          ��       ���   �        "�          ŀ       #�          #`       ���   72�       ܐ         ��        �          <�\       ��p   H�`       #�          �ǀ      ��          ?��       ��   ?r�        �          !        �          ! @       �    H��       �h           �      �           �       �   wy@        H            �      ��          �,        �   H��       ��           �      �          ��       ��   y         @            �      �                    �   ��       ��           `                    X        `   7|�       �0            @                             @   ��        �           �                    x        �   ?|�                     @                             @   �`       ��            �        �           ,         �   7~@       ߐ                                              (��       
 �            �        �           <         �   |@       
 �                                              '�       #l            P        �                    X   ?~        H                     �                       ?��       ��            p        �                    x                                  �                       �P       �                     @                    ,   x       �                      @                       �p       �                     �                    <            �                      @                                                         �                                                                                                                    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       ��  �    |�          �      �           ��  �    |�                                                                                                                                                                                           �  ` �    ��          `      l           �  ` �    ��                                                                                                                                                                                           �  ` �    ��          `                 �  ` �    ��                                                                                                                                                                                           �y�s��    ���?�       g��<|    ����       �y�s��    ���?�                                                                                                                                                                                        ��fl�    �홶ـ      �۶f�    ٛm�       ��fl�    �홶ـ                                                                                                                                                                                       �}�g��    �͙�߀      �6~�    ٛm�       �}�g��    �͙�߀                                                                                                                                                                                       �ͳf�    �͙��       �6`�    ٛm�       �ͳf�    �͙��                                                                                                                                                                                        �ͳfl�    �͙�ـ      �6f�    lٛm�       �ͳfl�    �͙�ـ                                                                                                                                                                                       �}�3��    |͏6�       �3<|    ���l�       �}�3��    |͏6�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �              �                           �              ��              �                           �              �                                                                                                                          �              �                           �              ��              �                           �              �                                                                                                                          �              �                           �              ��              �                           �              �                                                                                                                          �              �                           �              ��              �                           �              �                        � ��                 x 0 x                                                                   �              �                           �              ��              �                           �              �     3` <                 6 �0                 ̀0 �                                                                   �              �                           �              ��              �                           �              �     0`                   � 0                 ��0                                                                    �              �                           �              ��              �                           �              �     0sl�                 6� 0                 �ͳ�                                                                   �              �                           �              ��              �                           �              �     cm�                 �6ـ`                 y��`8                                                                   �����     �����      ����      ����       �����     ����������     �����      ����      ����       �����     �����     cm�                  66߀�                 ���                                                                                                                                                                                                  cm�                  66��                 ��                                                                                                                                                                                                   3a͘                 6ك                  ͇6`�                                                                                                                                                                                                  1��                 ���                 x�3�x                                                                                                                                                                                                   �                                                                                                                                                                                                                                                                      p                                                                                           