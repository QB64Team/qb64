��Z  �  ���>��00��>  ��@@��  ����  ���  �    ���   �� � ���G��6��?������?�������>��  �����        ���>��00��>"�"����EDED����ğ��"�2������  @��   �� � ���G��6��?������?�������>��  �����        ���>��00��>  ��AED���FG�Gď������������PP���
��#����h.�<���2r���8<|x���>�?�������>��  �����        ���>��00����  ����@@����@@�����������~�����}|�~������ ����@ ���� @����  ���� 0 ����� ����              ������� � �����  ������ � ���x��� @ @������      ������@ @ ������@ @ ������� � �����������������  ���������������   ���������   ���� � ������ � �����@ @ ������@ @ ������      ������ @ @������ � ���x���  ������� � ����������>�>�>�>        ������� � �����  ������ � ���x��� � �������   �������@p@������@�@п�(����	����p�����������&�>������L�|���������������0��������`�������D�G��?����I�O������;  ?  ������ @ @������ � ���x���  ������� � �����               p  p ������� � �3����S s ������P�p���x���P@p@￸��� P  p ߿����@P@p������@P@p�������P�p������P�p������P�p������P�p������P�p������P�p������P�p�����@P@p������@P@p������ P  p ߿����P@p@￸���P�p���x���s s ������� � �����                    ������� � �����  ������ � ���x��� @8 @������$  <  ������r ~ ������Y _ ����������s������@��y������ ��|���������~��������?�����d�|������2�>�����@@������@�@������� � ����������8�������x���  ������� � �����                                                                          ����            ����           ����            ����            ����            ����           ����            ����            ����            ����            ����            ����           ����            ����            ����            ����            ����            ���� (   <      ���� >         �_� ߀  ��     ��� �  ��     ���� ��  ��     �e� c   ��    ��?���  � ��               ����            ����           ����            ����            ����            ����           ����            ����            ����            ����            ����            ����           ���� (   <      ���� >         �_� ߀  ��     ��� �  ��     ���� ��  ��     ��    ��     �A� ��  ��     ����          ���� "   >      ����            ���� c        ��?���  � ��               ����            ����           ����            ����            ����            ����           ����            ����            ����            ����            ���� >          ����   ?     ���� ߀  �   �  ���� ��        ������      ���� ��        ���� ��        ���� Q   ?     ���� >        ����            ����            ����            ���� c        ��?���  � ��               ����            ����           ����            ����            ����            ����           ����         ���� 	   	   	  ���� �   �   �  ���� @  @  @ ���� ~   @   @  ����   	   	  ���� ��  ��  �� ����׀ >�  � ����� ?  ����߸ ?8 8 ���� ��  <@  $@ ����    A   A  ���� ��  ��  �� ����            ����            ����            ���� c        ��?���  � ��               ����            ����           ����            ����            ����            ����           ����         ���� Y          ���� ��         ����@         ����	~          ����         �����   �   � ������         ������         �������        ������         ����
         ���� ��         ����           ���� ��         ����"         ���� c        ��?���  � ��               ����  @   @   @ ����           ����            ����            ����            ����           ����         ����(Y          ����D��         ���� @       ����I: �        ����0E         ������   �   � �����@   @   @���� �         ���� ��        �����          �����  �   �   ���� ��         ����           ���� ��         ����"         ���� c        ��?���  � ��               ����            ����           ����            ����            ����            ����           ����            ���� @          ����@�          ����            ����@           ����           �����          ����            ����          ����  (         �����          ����          ���� ��         ����            ����  �         ���� "         ���� c        ��?���  � ��               ����            ����           ����            ����            ����            ����           ����            ����            ����            ����            ����            ����           ����            ����            ����            ����            ����            ����            ����            ����            ����            ����            ���� c        ��?���  � ��                                                                                                                                                                                                                                                                                                                                                                                                                             