��g  ��Q Q  g�����0   �    �                         �������   @ ?�                        ����d   ��� �      ?�                 n��?���    ?� D    ��                �������   c���                      ���  <���  H����	     ` �               _�p  /�`  �|  0�  � �@�             ���  ���  @�  �   �@0 @            ��    q��  g�   �    ���� �            �\    ��  �    = P    ���              ��    �� �    �   C���a             /�`    ?� p      �������             [��    �� $�    �  �A���              ��      ���(	�    �
 @ �B���0            ��      w��@      �  �B�             o�      ;� �&      8�  �B� �            _�      7� �l      6� �`��
�            ��      �� X      ; @ �P��            ��      ��@�      �  @`(��
            ~       ?��0      @  �0(��(4�            @  `  ���`  p  �  �($��HH�          � ��  �
  ��  �
�    t�� �           ��  ��  ��  ��� `  
p �     p   @ �      ���  ��� � `	
p$@<`           �        ���  �  � 8�� X��`            �   �L�  ׀   泀 � H��`0     �@�   �  ���  _�  �3�  � �$���0     ���   �  � �  k�  ���  � A  d�       @   �  ���  +�  ���  l ��� �     � �   �  � �  /�  ���  l  LO��0     � �   �  ��� ��  �� �  #_���@     � �   �  ������,  �!���  �=��       |   �  ?�~ 7�,  ?� � 6 �~�?�     >  >   �  >�> ��,  ? ~ �6 o|�ߟ      <     �  z@�/ �\  z�b� ;  �}^�_      x     �  ���� �X  ��P� ;  z��       �    �  ��  �X       �����          �  ���| �X  X|    0�����           �  s���X  ��   �_�w�      �    �  (�
 ˀX  " �   �����           �  X����X  "�� '�������           �  (�
  �X  "   '� �����           �  S�` �X  �`   ? �_�w�      �    �  �ǈ �X  	H    ������           �  �� �X      ����           �  ������X  �P��   z��             �  zs��8�  z���8   �}\_      x O   �  >�.`��,  > .`�4  }���      <     �  ?�~��,  ?  ~� ������      >  >   �  ������,  � ��� � �}�~        |   �  ���D �  �c�D 4  ���      � �   �  7��� +�  7��� (  ���      ��   � ������/� ������l  0��      ��   � ���C@/� ���C@h  @���      ���   � �!��� �W� �!�� �P   ���  8     ��   ��F���x_��F���x�   �   0     >�    � ��Đ��� �tĐ�   �   p     p     �82)��H���2)��H�         `            ��BR��$_��BR��$@         �          @ ������� �����`         �          @ `��J
���`��J
�  �      �          � p	�I���p	�I�  �      �         � ��8
$�E���@�8
$�E��  `                  ��`(�E��� L`(�E�  0                  ���((�B���� 6�((�B��                    ���(P�A�o�� �(P�A�l                    �� PP�A@_���PP�A@�        (           ���`P������@�`P����        p         0  �`�`����  `�`���`   �     �         `  =������f�� �����f�   �    �   �     �  �ɀ���)�  ̀���)    p    �    @       �� ��`7��   w ��`7     8         0       ����`��x  �9���`� �       <            ��a��c7��  q��c4 @   �   �         0   �����|���  ���|�    �  �     �   �   ��c���_��   c���`      �  �      `       ���?���    \?��     ?��              }������    ��       ���       ��     �������      ���        �         ?�      �������   @ �                          �������                                                                   Q Q  g�����0   �    �                         �������   @                           �����d   �     �                         n�������         D                        �������    �                         ��������  H �� 	      �                _�����`  � � �   ��              ��������  @ q���       8  @            ���  8���  ����    � p �  �            ��p  ?��  ~  ?  P   �����              ���   ���  �  �     ���`             /��    g��  �  �    ���              [��    �� $ g    r    ����              ��X    ���( �     
 @  ��� �             ���    ���@�    
�  @`���             o�@    ?� �p     � �`�� �             _��     �� ��    ��  P�� @             ��      _�� �     � @@0��
              ��      _��@      X   `(b�0           �      O���      L   0(R�8            �  `  %���&  p  &   �((            ��  �
  �� l  �
�    r�H�           ��  ��  �� X  ���     
p       p    �     	� �  ��� 	�  `	p"@           ��      �� �  �  �  L�  ,�{            �@  �L� ��P  泀 �  �H����     �@�  � �@ ��� ��` �3� �  ��$����     ���  � �@ � � ��` ��� �  ���  ds�      @  � �� ��� _�� ��� `  XO� �� �    � �  @ �� � � �� ��� `  &/�� �    � �  @ �� ��� /� � �� 0  ?���` �    � �    �  ��� ��� �!� �  �=�� `      |    �  ?�~￀� ?� �� `>�>0 `    >  >    �  >�> �� ? ~ � ~|�ߟ� `    <      �  z@�/ ��� z�b� � ��^�_  `    x      �  ���� W�  ��P� X �z��  0     �    �  ��  W�    X  a���� 0         �  ���  _�  X  X  ����� 0          �  s� _�  � X  �_�w� 0     �    �  (�
 �_�  " �X   ����� 0          �  X��߀  "�� ������� 0          �  (�
  [�  "  \ � ����� 0          �  S�` [�  �` \ ��_�w� 0     �    �  �ǈ [�  	H \  ����� 0          �  �� _�   X  ���� 0          �  �����_�  �P��X  z��  0           �  zs��0��� z���0� �}\_  p    x O    �  >�.@���� > .@�� ?����  p    <      �  ?�~ ��� ?  ~ � �~���  `    >  >    �  ��� ��� � � �  �}�~  `      |    �� ����/�� �c��0  ���  �    � �    �� 7��&_�� 7��&@  ���  �    ��  @ ��������������`  0��  �    ��  @ �@��Ԇ���`��Ԇ��  ����� �    ���  � �@p&���AB��`p&��AB�  �  ��� �     ��  � �c�I?�I 俀s�I>�I ��  �  �  �     >�   � �� �7�H�5�� �7uH�5   @  �  �     p    ��bJ�$P	�� �bJ�$P	�  @                  �X�R��(
� ��R��(
�                     ������� L���   0                  �	��
&���&	��
'                     �
��i���3
��j                     ��(��W��@�(��T         8           ���((����� 
�((���        p            ��@00��_�� @00��P   �     �         @  ���P0������ �P0����   �    �    �     �  ��X`P�����X`P���@   �    �    @       ��$�`�@����@ ��`�@��   x                 ���`�����   S�`���     <                =���@�����  �@���         |            ��p���'��  
p���$    �   �             ���������   �����     �  �     �   �   �q���_�x  � q���` �    �  ?�      p      �������   ,�  @    ��             ��������   ��      ���       ��    ���������    ���        �         �      ���������     �                           }�������                                   �������                                    �������   @                             �������                                                                   Q Q  g�����0   �8  �                         �?���}�   @�  �                      ~�����d   �    @�                        n������       D                        ��������                            ���������  H@    	                        ^������`  �  �  B�  �     �             ���`���  B  �� !     �   @            ����/���   �0     � �� �            ���������  1��� P      8               ��O� ���  ����    0 �             /��8  ��  ?  >    �����              [���  ��� $@�  �    ���`              ���@   ����( 	�  � 
 @� ���0 �            ���    7���A     t A  `���             m��    �� � N    9 $�  0 ��              _�8    � � �    �� @0��              ��0    ?�0    @ @ �(��
�             ��`    ��H`       ����            ��    /����    0  b��            o�� ` ����� p �   �(8`             ��  �
  ���� �
� �   
r�PPp           ��  ��  K��   ��� �  
p�8      p    ��     +��   ��� h   p"@           ��      7��@,  �  6   �  $�            ��  �L� ��@,  泀    D�� n      �@�   � ��� ���X �3�  @#�����      ���   � � � 
���X ���     ��  d�       @   � ��� ��0 ��� �  @PO� ��     � �   �  � � �� � ��� �  @,/��     � �   �� ��� � � ��    @���`�    � �   �@ ��� >�� ` �!� >�  ��=���      |  � �` ?�~���` ?� ���  �>�>p�    >  >  � �@ >�>���` ? ~��  �|�ߟ��    <    � �@ z@�/��` z�b��  ���^�_ �    x    � �� ����_� � ��P�`  �z��  �     �   @ �� �� ��  `  0���� �        @ �� ��� �� X `  ����� �         @ �� s�|�� �|`  �_�w� �     �   @ �� (�
��� "�`   ����� �         @ �� X���� "�` ?������ �         @ �� (�
 o�� " p ? ����� �         @ �� S�@o�� �@p  ��_�w� �     �   @ �� �ǈ0�� 	H0`  ����� �         @ �� ���� `   ���� �         @ �� ����_� � �P�`  z��  �          @ �@ zs��¿�` z���  ��}\_ �    x O  � �@ >�.����` > .���  ����� �    <    � �` ?�~`>��` ?  ~`>�  ��~��� �    >  >  � �@ ����� ` � ��  ��}�~ �      |  � �� /����� � /�c��   @��� �    � �   � ���4�� ����4�  @���      ��   ������0����  @`��      ��   �8��Ć����X8��Ć�    ����      ���   ��$���A����X�$��A� @#  ���       ��   �� I?�Q t��@. I>�Q u     �        >�    �� �7�H���@. �7uH�     �        p    ��BR��P/�� BR��P,                     ������(K�� ����(L        8            �������	����         8            o������������         p             w�X
(��_���X
(��@  �     �         @  �� (����@0(��@   �    �         @  ���0�����  �0���   �    �    �     �  ���00��߀ L00���    p         @       ��� `��6���  6 `��7     8         0       ���``��I��� 	�`���        <            ���`����}�@��`�Ü �       p            ��0���o��   8���p     �  �         `   =���������  �����      �  �      �  �   ���������  ���ƀ    ~  ?       0      ����;���    n�:       ��         8    {������x  � �� �    ���       ��    ���������   ���  @     �         �     ������{�  � �  �                        ���������                                   ���������                                }�������                                   �������                                   �������   @                            �������                                                                   Q Q  g�����0   �8  �                         �?���}�   @�  �                      ~�����d   �    @�                        n������       D                        ��������                            ���������  H@    	                        ^�������`  �      B�  �     �             ���������  B      !          @            ���������            �      �            ��������   �  P                       ��������  ��      �              /����?���   �0    ��               [�������� $@ ���       0               ����  1���(  G�� 
 @� 8 �  �            ����  ����A �  <� A   `@�              m��`  ?�� � x  0 $�  �A� �              _���   ��� � �  � �  a� `              ���    o�� �   �  @ 0a�              ���    ���H     v    a�             ��    ���� .    ;    a�             o�� ` ���� X p �     �              ��� �
  ��� � �
��    Dr�03             ��@ �� _�� P ���`   �pP�      p    ��@    ��� ` ����   �p!A�         �  ���    ��@� � p   �  B��          @  ��  �L� ���@� 泀�    � `      �@�    � ��� ����	��3� � @ ���p      ���    � � � S��� ��� �   �S  d8       @   � ��� S��� ��� T   p/� �|8     � �   �� � � /��  ��� l   ���     � �   �� ��� +��  �� (   ���@     � �   �� ��� ��  �!� 6   �=��       |   �� ?�~��� , ?� ��   ~�>      >  >   �� >�>?��� , ? ~?�    ��ߟ�     <     �� z@�/�� , z�b�   �}^�_      x     �� ����
�� X ��P�    �z��       �    �� �� 
�� X      ����          �� ��� 
�� X X     �����           �� s�p�� X �p    �_�w�      �    �� (�
��� X "�     �����           �� X���� X "�   '������           �� (�
 �� X "    '������           �� S� � X � �   ?�_�w�      �    �� �ǈ`�� X 	H`     �����           �� ��
�� X     ����           �� ����
�� X �P�    z��             �� zs����� , z����   ��\_      x O   �� >�.���� , > .��   �}���      <     �� ?�~@�� , ?  ~@6    ~���      >  >   �� ������  � ��4    �}�~        |   �� o���P+��  o�c�P(   ���      � �   �����</�� ���<l   ���      ��   ����S������T   0�� 8     ��   �0���_���0����   @��� 0     ���   �@(���������(���� @  ��� p      ��   ���P��Q@���@�P��QA�     �  `      >�     ����W�P�O��@��WuP�P     �  �      p  @  ��a���(b�� q���(b`   �    �          @  ��3��6��� 3��6�   �    �          �  ����������    `         @       o�(���� ���    p                 w��(�6���� W(�7    8                ���0�m���@ +�0�n                     ���0������  �0���        p            ���p0��7�߀ 
p0��8     �   �             ����`������  �`���     �  �     �   �   ���F`��?��� G`��@     �  �      @      ��y����}�@� ���΀ �    >  ?       8      ����1���    ~�2       ��         0    =��������   ��       ���       ��    ��������   ��`      ?��        �     ��������     ?��                          {�������x  �      �                       ���������         @                       ������{�  �     �                        ���������                                   ���������                                }�������                                   �������                                   �������   @                            �������                                                                   Q Q  g�����0   �8  �                         �?���}�   @�  �                      ~�����d   �    @�                        n������       D                        ��������                            ���������  H@    	                        ^�������`  �      B�  �     �             ���������  B      !          @            ���������            �      �            ���������       P                       ���������                            /���������                              [��������� $@  �                         �����?����(  ��  
 @�  �   �            �����o����A  �p  A    ��              m�������� �  8���  $�     p               _��g� ���� �  ���  �   �               ����  �� �  }�  @    �               ���0  ���H <  @     � ��             ��@  ����� p  �    �1� @             o���` ����� �p�     �               ��� �
 o��� ��
��     q�             ��� �� ���   ���T    
p0(       p     ���   3���  . ���2     pP�             ���    ���@ L �      1�  ��             ��� �L�
���@ X 泀
      �       �@�   ��������� ��3�� @ @b��       ���   �@� �����P����    �S  d�       @ �  �@�������`����    �/� �=�     � � �  ���� ���  ����@   ����     � � @  �������� ���`   ���`�     � � @  ������_�� ��!�@   �=���       | @  ���?�~��� �?� ��   ��> `     >  >    �� >�>��� �? ~�    |�ߟ p     <      �� z@�/��� �z�b��   `}^�_ p     x      �� ������� ���P��   ~z�� 0      �    �� �� ���   �   ����0          �� ��� ���  X �   �����0           �� s� ���  � �   �_�w�0      �    �� (�
|_��  "|X    �����0           �� X����  "�   ������8           �� (�
 W��  " P   ������8           �� S� _��  � X   �_�w�0      �    �� �ǈ ���  	H`�    �����0           �� �����  �   ����0           �� ��ж��� ��P��   z�� 0            �� zs����� �z����   �\_ p     x O    ���>�.��� �> .�    }��� `     <      ���?�~��� �?  ~��    ~��� `     >  >    ������A_�� �� �A@   �}�~ �       | @  ���������� ���c��`   ��� �     � � @  �����s��  ���s@   ��� �     �� @  �H�������h����    ����     �� �  �`�������p����    �����     ��� �  ��(������ �(�⍀ @ @ ���       ��   ��Xq?�!����@ �q>�a��      �        >�    ������P����@ L��vP�     0 �        p    ��炊�0w���  '���0v                      ����(o���  ;�(l                    �������� ���         0            o��L�	?���� L�	0     �   �             w��8����� 8�`    �  �         @   ����0�����@ �0��      �  �      �  �   ����0�r����   �0�r�     x                �����Ǐ��߀  x�ǎ         |             �����w����   �t       ��         p    ����������  ��      ���        ��    ��������}�@� ���  �     ?�         �     ���������     �                           =���������                                 ���������                               ���������                                  {�������x  �      �                       ���������         @                       ������{�  �     �                        ���������                                   ���������                                }�������                                   �������                                   �������   @                            �������                                                                   Q Q  g�����0   �8  �                         �?���}�   @�  �                      ~�����d   �    @�                        n������       D                        ��������                            ���������  H@    	                        ^�������`  �      B�  �     �             ���������  B      !          @            ���������            �      �            ���������       P                       ���������                            /���������                              [��������� $@                             �����������(        
 @�       �            �����������A        A                     m�������� �   �   $�                      _������� �   p�  �   �                �����o���  �p   @   ��               ����������H  ���        `              ���  g�����  pf       �              o���`�����  o��        �               ����
����  ��
��      `q�              ���`�����  x���@     �p0�       p     ���� ����  ����     p`@             ���    _���@ @�P     �  ��              ��� �L�����@ �泀�     A��P       �@�    �����W���� �3�T  @ `��8       ���   ��� �)���� ���*     3  t        @   �����7���� 
���6     � �      � �   ���� ����  ,���     ��n      � �   ���������  X��     &����      � �   ������
���  X�!�
     #�=��        |   ���?�~��  (?� ��    @��>      >  >   �� >�>���  �? ~�    @|�ߟ      <     ���z@�/���  �z�b��     @}^�_�     x     �������?��  ���P�@    Lz���      �    ��@����� `�    ����        �  ��@������ `X�    �������         �  ��@s���� `��    ��_�w��      �  �  ��@(�
r��� `"r�    �������         �  ��@X�~��� `"~�    �������         �  ��@(�
��� `"�    �������         �  ��@S���� `��    ��_�w��      �  �  ��@�ǈB��� `	HB�    �������         �  ��@��2��� `2�    ����         �  �������?��  ��P�@    Oz���            ���zs����  �z���     @}\_�     x O   �� >�.���  �> .�    @}���      <     ���?�~���  (?  ~��    @~���      >  >   ����������  X� ��     !�}�~        |   �������k���  X��c�k     #���      � �   �����4���  .��5     ���      ��   �����'���� *���&     ��      ��   �����/���� ���,     ���      ���   ��0���s���� 0��t  @  ���       ��   �����a����@ ྾a�      � 0       >�    ������a����@ ��va�      � `      p     ���!�2���  !�2`     �  �         @   ���������  ���     �  �      �   �   ���������  ���      x         `      o��Ә�������  S���       <               w���p������  <p�      � �             �����k����@  �l       ��         `    ����������   ��      ���        ��    ����O���߀   ���        ?�         �     �����������    �                           �����������                               ��������}�@�       �                       ���������                                  =���������                                 ���������                               ���������                                  {�������x  �      �                       ���������         @                       ������{�  �     �                        ���������                                   ���������                                }�������                                   �������                                   �������   @                            �������                                                                   Q Q    <�       � �       @                  �đ�      ;n        �                 >�>`      �� ��      @                  �����               @                ;��f     �l�      �                 L�?�_�     3��f      � @�               �������    @       �  �              g�����`    �   �     @                  ����?�   �   �`                        ;�����h   �    �                       �������                @              =�������                               [�������   $  ?�    @                  ��`?�v�  H��� �      �                n���o��@  � �p D�  @  ��              }������`  � ���  �  !   p B             ��'  p�� D ��� @    �               ���  �� @�  }�      �              ��0  _�� <  `  � � �� �            
���  ���  �  � P 1� @             ���` ��� 	 �p�@  �              �� �
 k�� 
@��
��    q�             +�� �� ��  5 ���T    @
p0(      p     ;�   3�� �. ���2   pP�             W�    �� (�\ �    !�  ��              W�P �L�
� ( � 泀
�@   �       �@�   ��������	 ��3�  @ @b���      ���   ��@� ����BP����  �S  d�       @ �  ��@����߀P`����   �/� �=�     � � �  ���� �_� R����` ������     � � @  {�����_������@  ���`�     � � @  _�����_��!�@ �=���       | @  [��?�~ �����?� � �   ��> `     >  >    �� >�>�� �? ~��� |�ߟ p     <      �� z@�/��@�z�b�� `}^�_ p     x      �� �������H���P��   ~z�� 0      �    �� �� W��H  X   ����0          �� ��� _��  X X	 H�����0           �� s� _��H � X   �_�w�0      �    �� (�
|_��H "|X    �����0           �� X����  "�	 H������0           �� (�
 _��H " X   ������0           �� S� _��H � X   �_�w�0      �    �� �ǈ _��  	H`X	 H �����0           �� ��_��H X   ����0           �� ��ж���H��P��   z�� 0            �� zs����@�z���� �\_ p     x O    �� >�. �� �> . ��� }��� p     <      [��?�~ �����?  ~��    ~��� `     >  >    _�����AO�� �AP �}�~ �       | @  {�������������c��`  ��� �     � � @  �����s_� R ���s` ����� �     �� @  ��H����߀Ph����   ����     �� �  ��`������Bp����  �����     ��� �  ���(�������	 �(���� @ @ ���       ��   W�Xq?���� ( �q>�a� @    �        >�    W����P��� (�\��vP�     �        p    ;ǂ��0w�� �'���0v                    +���(o�� @�(l                    ������� 
 ���         0            ��L�	���  L�	�     �   `             �������  ���   @   @         @   ��0���x  ��0�� �    �  �      �  �   ���0�r���   �0�r�     x                ����ǎ���   X�Ǐ       ?  |             ����u���  ! 7�v B     ��         p    ��������  @ ��      ���        ��     ���������    ���        �         �      w�������   @ �                          /�������                                �������         @                         �������                                  �������                                   �������     @                             w�����@    �  �                          ~���      � @�                           /��o��      �                            �����       @                           �����      @                              ��o��       �                             ;���       @                                                          Q Q    <�       � �       @                  �đ�      ;n        �                 >�>`      �� ��      @                  �����               @                ;��f     �l�      �                 L�?�_�     3��f      � @�               �������    @       �  �              g�����`    �   �     @                  ����?�   �   �`                        ;�����h   �    �                       �������                @              =�������                               [�������   $        @                  ������v�  H�     �                        n������@  �  �  D�  @                   }��0��`  �  ��  �  !  �  B             ����o�� D �p @    ��               �������� @ ���       `              ��Ӏ ����  3��   �  �  �            
��N  9��   �  y� P  0�              ���`��� 	 �p�@   @ �              ��`�
_�� 
@p�
�`     �q��             +��������  �����    @p0`      p     ;��  ��� ������   p`              W�    o�� (� � h   �� ��              W�� �L�g�� ( 7 泀d @  A��       �@�    ������3���	 .�3�2  @ `��       ���    ���� ����B L���   03  t        @   �������߀P X���     � �      � �   ��P� �
�� R ����
  �� $��7      � �   {��������� ����   G����      � �   _����� ��!�   C�=�~��       |   [�`?�~����`?� ��    ���?�     >  > �  ��@>�>�� `? ~��� �|�ߟ�     <   �  ��@z@�/~��@`z�b�~�  �}^�_�     x   �  ��@�������H`��P��    �z���      �  �  �����_��H�`   �����        @  �������� �X`	 H������         @  ���s���H��`    �_�w��      �  @  ���(�
s��H�"s`    ������         @  ���X�_�� �"@	 H?������         @  ���(�
_��H�"@   ?������         @  ���S���H��`    �_�w��      �  @  ����ǈA�� �	HA`	 H ������         @  �����;��H �;@   �����         @  ��@�������H`�P��    �z���          �  ��@zs����@`z����  �}\_�     x O �  ��@>�.��  `> .��� �}����     <   �  [�`?������ `?  ��    ������     >  > �  _�����E �� �E   A}�~�       |   {�0�������� ���c��   G���      � �   �����:�� R X��:  �� $���      ��   �������߀P X���     ��      ��   ���������B ,���   ���      ���   ���0���%���	 .0��&  @  ���       ��   W��a?����� ( a>��� @   �        >�    W����`��� (���t`�    � 8      p    ;���!��� �
��!�       p             +��c�3O�� @c�3P    �   �         @   ������� 
 ���     �  �      �   �   ��L�?��  L�@      �  �      @      ��3�����   ����    |         0      ���ϙ��x  � ,�Ϛ  �      |             ����g���   �h      ��         `    ���p���   p        ���        p     ���������  !  O�  B      ?�         �     ���������  @  �                           ���������                                   w�������   @                             /�������                                �������         @                         �������                                  �������                                   �������     @                             w�����@    �  �                          ~���      � @�                           /��o��      �                            �����       @                           �����      @                              ��o��       �                             ;���       @                                                          Q Q    <�       � �       @                  �đ�      ;n        �                 >�>`      �� ��      @                  �����               @                ;��f     �l�      �                 L�?�_�     3��f      � @�               �������    @       �  �              g�����`    �   �     @                  ����?�   �   �`                        ;�����h   �    �                       �������                @              =�������                               [�������   $        @                  ������v�  H�     �                        n�������@  �      D�  @                   }�������`  �       �  !      B             �������� D      @                      ���0��� @  ��      �               ����_���  �`   �  ��  �            
��������   ���  P    `              ��Ӏ ���� 	  3�� @    �              ��� 
��� 
@ o�
�      p�              +��X����   �����    @  p       p     ;�  ?�� �(���@    �p!�             W�@  �� (�p�    �  `�              W����L���� ( �況� @  ��`       �@�    ����������	 ��3��  @  ��p       ���    ���� �����B 
�����   3  t0        @   ������K�߀P ���L    � �8      � �   ���� �+�� R ���(  �� ��      � �   {�����5���� *��6    ����      � �   _������ ,�!�   �=��        |   [��?�~���� \?� �      ��>      >  >   ���>�>
��  X? ~ ��  |�ߟ      <     ���z@�/���@ Xz�b��    }^�_      x     ��Є������H X��P�     &z��       �    �� ����H ��    G����           �� �����  �X�	 H @�����            ���s����H ���    @�_�w�       �    ���(�
e���H �"e�    @�����            ���X�}���  �"}�	 H O�����            ���(�
���H �"�    O�����            ���S����H ���    @�_�w�       �    �� �ǈ��  �	H�	 H @�����            ��0��M��H �M�    A����            ��X������H ؅P��    'z��             ���zs����@ Xz���    }\_      x O   ���>�.��  X> . ��  }���      <     [��?����� \?        ~���      >  >   _������� ,� ��   �}�~        |   {���������� .�c��    ���      � �   �����)�� R ��j  �� ���      ��   ������O�߀P ���L    ��8     ��   ����������B �����   ���8     ���   ������ï���	 ��è  @  ���p      ��    W��A?�AW�� ( a>�AX @  �� �      >� @   W�1��fo�� (�1�vfp   ���      p @   ;���-��� ���-�    �  �      �  �   +����2��� @��2�     x                ��S����� 
  ����      <               ���p����   lx�       � �             ����k���   �l     ��         `    ������x  � ��  �    ���        ��    ���������   ���       ?�         �     ���������    ?�                           ���������  !      B                        ���������  @                               ���������                                   w�������   @                             /�������                                �������         @                         �������                                  �������                                   �������     @                             w�����@    �  �                          ~���      � @�                           /��o��      �                            �����       @                           �����      @                              ��o��       �                             ;���       @                                                          Q Q    <�       � �       @                  �đ�      ;n        �                 >�>`      �� ��      @                  �����               @                ;��f     �l�      �                 L�?�_�     3��f      � @�               �������    @       �  �              g�����`    �   �     @                  ����?�   �   �`                        ;�����h   �    �                       �������                @              =�������                               [�������   $        @                  ������v�  H�     �                        n�������@  �      D�  @                   }�������`  �       �  !      B             �������� D      @                      ��������� @                            ��������   �    �       �            
��������    p   P   �               ��������� 	  ��� @    p               ���p/��� 
@ �0      � �               +���������   ���     @   0              ;�� u��� � 7���     p              W��  ��� (� N�9     1                 W��0�L��� (  �泜� @   A��        �@�    ���a���?���	 q�3�@  @  ����       ���    ���A� ß���B a��à    �  l�        @�   �������_�߀P ����@    � ��      � �@   ����� ���� R Ͽ���  �� ��`      � �    {���������� ����    ���p      � �    _�����_� �!�X   �=��        |   [��?�~W���� ?� �P     ~�>8      >  >   ���>�>o��  ? ~h �� |�ߟ      <     ���z@�//��@ z�b�,   }^�_      x     ���������H ��P�     z��       �    �����7���H 4     ����           ���������  ,X 	 H �����            ���s����H ,�     �_�w�       �    ���(�
���H ,"     �����            ���X�w���  ,"v 	 H �����            ���(�
���H ,"     �����            ���S����H ,�     �_�w�       �    ����ǈ5���  ,	H6 	 H �����            �����u���H ,v     ����            ���������H �P�     	z��             ���zs��+��@ z���(   }\_      x O   ���>�.k��  > .l �� }���      <     [��?�~W���� ?  ~P     ~���8      >  >   _������� � ��   �}�~0        |   {���������� ��c��    ���p      � �    ��������� R ����  �� ���`      ��    ���O���_�߀P O���@    ����      ��@   ���9��Ɵ���B 9��Ơ    �����      ����   ������̿���	 ����  @  �����      ����   W��M��Y�� (  ;�Y� @   p�       @>�    W���f��� (� wtg     8�       0p    ;�Ɉ����� � )���       <             +���x�3��� @ x�4      � �         0    ��������� 
  ���       ��       � �    ���p?���   p@        ���        p     ���������    O�       ?�         �     �������x  �  �   �                       ���������                                ���������                                 ���������  !      B                        ���������  @                               ���������                                   w�������   @                             /�������                                �������         @                         �������                                  �������                                   �������     @                             w�����@    �  �                          ~���      � @�                           /��o��      �                            �����       @                           �����      @                              ��o��       �                             ;���       @                                                          