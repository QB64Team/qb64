��   �                                                                                  ����������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                      ���������������������������������������������������������������������������  �����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������   �����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������   �����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      �������������������������������������������������������������������������     ����������������������������������������������������������������������������                                                                                                                                                                      �������������������������������������������������������������������������      ���������������������������������������������������������������������������                                                                                                                                                                      �������������������������������������������������������������������������      ���������������������������������������������������������������������������                                                                                                                                                                      ������������������������������������������������������������������������       ���������������������������������������������������������������������������                                                                                                                                                                      ������������������������������������������������������������������������        ��������������������������������������������������������������������������                                                                                                                                                                      ������������������������������������������������������������������������        ��������������������������������������������������������������������������                                                                                                                                                                      �����������������������������������������������������������������������         ��������������������������������������������������������������������������                                                                                                                                                                      �����������������������������������������������������������������������         ��������������������������������������������������������������������������                                                                                                                                                                      �����������������������������������������������������������������������          �������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������           �������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������           �������������������������������������������������������������������������                                                                                                                                                                      ���������������������������������������������������������������������             ������������������������������������������������������������������������                                                                                                                                                                      ���������������������������������������������������������������������             ������������������������������������������������������������������������                                                                                                                                                                      ���������������������������������������������������������������������             ������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������               ��������������� �������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������               ��������������   ������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������� �������������                 ������������    ������������������������������������������������������                                                                                                                                                                      �����������������������������������������������������  ������������                 �����������     ������������������������������������������������������                                                                                                                                                                      �����������������������������������������������������   �����������                 ���������       ������������������������������������������������������                                                                                                                                                                      �����������������������������������������������������    ���������                   �������       �������������������������������������������������������                                                                                                                                                                      �����������������������������������������������������     ��������                    �����        �������������������������������������������������������                                                                                                                                                                      �����������������������������������������������������      ������                      ���         �������������������������������������������������������                                                                                                                                                                      ������������������������������������������������������      �����                                  �������������������������������������������������������                                                                                                                                                                      ������������������������������������������������������                                             �������������������������������������������������������                                                                                                                                                                      ������������������������������������������������������                                             �������������������������������������������������������                                                                                                                                                                      ������������������������������������������������������                                             �������������������������������������������������������                                                                                                                                                                      ������������������������������������������������������                                            ��������������������������������������������������������                                                                                                                                                                      ������������������������������������������������������                                            ��������������������������������������������������������                                                                                                                                                                      �������������������������������������������������������                                           ��������������������������������������������������������                                                                                                                                                                      �������������������������������������������������������                                           ��������������������������������������������������������                                                                                                                                                                      �������������������������������������������������������                                           ��������������������������������������������������������                                                                                                                                                                      �������������������������������������������������������                                           ��������������������������������������������������������                                                                                                                                                                      �������������������������������������������������������                                           ��������������������������������������������������������                                                                                                                                                                      �������������������������������������������������������                                          ���������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������                                         ���������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������                                         ���������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������                                         ���������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������                                         ���������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������                                         ���������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������                                        ����������������������������������������������������������                                                                                                                                                                      ���������������������������������������� ����������������                                       ����������������������������������������������������������                                                                                                                                                                      ���������������������������������������   ���������������                                       ��������������  ������������������������������������������                                                                                                                                                                      ���������������������������������������   ���������������                                       ��������������  ������������������������������������������                                                                                                                                                                      ���������������������������������������    ��������������                                       �������������   ������������������������������������������                                                                                                                                                                      ���������������������������������������     �������������                                       ������������     �����������������������������������������                                                                                                                                                                      ��������������������������������������      �������������                                      �������������     �����������������������������������������                                                                                                                                                                      ��������������������������������������       ������������                                      ������������      �����������������������������������������                                                                                                                                                                      �������������������������������������         ������������                                     ������������       ����������������������������������������                                                                                                                                                                      �������������������������������������         ������������                                     �����������        ������������������  ��������������������                                                                                                                                                                      ����������������     ���������������           �����������                                     ����������         ����������������    ��������������������                                                                                                                                                                      ����������������            ��������            ����������                                     ���������           ������������       ��������������������                                                                                                                                                                      ����������������                 ��             ����������                                    ����������            ��������          ��������������������                                                                                                                                                                      �����������������                                ���������                                    ���������                              ���������������������                                                                                                                                                                      �����������������                                 ��������                                    ��������                               ���������������������                                                                                                                                                                      �����������������                                 ���������                                   �������                               ����������������������                                                                                                                                                                      �����������������                                  ��������                                   �������                               ����������������������                                                                                                                                                                      ������������������                                  �������                                   ������                                ����������������������                                                                                                                                                                      ������������������                                  �������                                   ������                                ����������������������                                                                                                                                                                      ������������������                                   ������                                   �����                                 ����������������������                                                                                                                                                                      �������������������                                  �������                                  ����                                  ����������������������                                                                                                                                                                      �������������������                                   �����                                  ����                                  �����������������������                                                                                                                                                                      �������������������                                    ����                                  ���                                   �����������������������                                                                                                                                                                      �������������������                                     �                                     ��                                   �����������������������                                                                                                                                                                      ��������������������                                                                                                               �����������������������                                                                                                                                                                      ��������������������                                                                                                               �����������������������                                                                                                                                                                      ��������������������                                                                                                              ������������������������                                                                                                                                                                      ���������������������                                                                                                             ������������������������                                                                                                                                                                      ���������������������                                                                                                             ������������������������                                                                                                                                                                      ���������������������                                                                                                             ������������������������                                                                                                                                                                      ����������������������                                                                                                           �������������������������                                                                                                                                                                      ����������������������                                                                                                           �������������������������                                                                                                                                                                      ����������������������                                                                                                           �������������������������                                                                                                                                                                      ����������������������                                                                                                           �������������������������                                                                                                                                                                      ����������������������                                                                                                            ������������������������                                                                                                                                                                      ����������������������                                                                                                            ������������������������                                                                                                                                                                      ���������������������                                                                                                             ������������������������                                                                                                                                                                      ���������������������                                                                                                              �����������������������                                                                                                                                                                      ��������������������                                                                                                               �����������������������                                                                                                                                                                      ������������������                                                                                                                  ����������������������                                                                                                                                                                      ������������������                                                                                                                    ��������������������                                                                                                                                                                      ���������������                                                                                                                          �����������������                                                                                                                                                                      ��������������                                                                                                                           �����������������                                                                                                                                                                      ��������������                                                                                                                           �����������������                                                                                                                                                                      ���������������                                                                                                                         ������������������                                                                                                                                                                      ����������������                                                                                                                       �������������������                                                                                                                                                                      �����������������                                                                                                                      �������������������                                                                                                                                                                      �����������������                                                                                                                    ���������������������                                                                                                                                                                      ������������������                                                                                                                   ���������������������                                                                                                                                                                      ��������������������                                                                                                               �����������������������                                                                                                                                                                      ��������������������                                                                                                               �����������������������                                                                                                                                                                      ���������������������                                                                                                             ������������������������                                                                                                                                                                      �����������������������                                                                                                          �������������������������                                                                                                                                                                      ������������������������                                                                                                        ��������������������������                                                                                                                                                                      ��������������������������                                                                                                     ���������������������������                                                                                                                                                                      ���������������������������                                                                                                   ����������������������������                                                                                                                                                                      ����������������������������                                                                                                 �����������������������������                                                                                                                                                                      ����������������������������                                                                                                ������������������������������                                                                                                                                                                      ������������������������������                                                                                             �������������������������������                                                                                                                                                                      ������������������������������                                                                                            ��������������������������������                                                                                                                                                                      �������������������������������                                                                                          ���������������������������������                                                                                                                                                                      ��������������������������������                                                                                        ����������������������������������                                                                                                                                                                      ����������������������������������                                                                                     �����������������������������������                                                                                                                                                                      ����������������������������������                                                                                     �����������������������������������                                                                                                                                                                      ������������������������������������                                                                                  ������������������������������������                                                                                                                                                                      �������������������������������������                                                                                �������������������������������������                                                                                                                                                                      ��������������������������������������                                                                              ��������������������������������������                                                                                                                                                                      ���������������������������������������                                                                            ���������������������������������������                                                                                                                                                                      ����������������������������������������                                                                          ����������������������������������������                                                                                                                                                                      �����������������������������������������                                                                        �����������������������������������������                                                                                                                                                                      ������������������������������������������                                                                      ������������������������������������������                                                                                                                                                                      �������������������������������������������                                                                    �������������������������������������������                                                                                                                                                                      ��������������������������������������������                                                                  ��������������������������������������������                                                                                                                                                                      ���������������������������������������������                                                                ���������������������������������������������                                                                                                                                                                      ���������������������������������������������                                                               ����������������������������������������������                                                                                                                                                                      ���������������������������������������������                                                              �����������������������������������������������                                                                                                                                                                      ����������������������������������������������                                                             �����������������������������������������������                                                                                                                                                                      ����������������������������������������������                                                            ������������������������������������������������                                                                                                                                                                      ����������������������������������������������                                                            ������������������������������������������������                                                                                                                                                                      ����������������������������������������������                                                            ������������������������������������������������                                                                                                                                                                      ����������������������������������������������                                                            ������������������������������������������������                                                                                                                                                                      ����������������������������������������������                                                            ������������������������������������������������                                                                                                                                                                      ���������������������������������������������                                                             ������������������������������������������������                                                                                                                                                                      ���������������������������������������������                                                              �����������������������������������������������                                                                                                                                                                      ���������������������������������������������                         ����                                 �����������������������������������������������                                                                                                                                                                      ��������������������������������������������                   �����������    ������                        ����������������������������������������������                                                                                                                                                                      ��������������������������������������������                ��������������    ����������                    ����������������������������������������������                                                                                                                                                                      ��������������������������������������������           �������������������    ���������������               ����������������������������������������������                                                                                                                                                                      �������������������������������������������     ��������������������������    ��������������������           ���������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    �������������������������      ���������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ������������������������������ ���������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ��������������������������������������������������������������������������    ����������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                      ����������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                    