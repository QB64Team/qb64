�i  $(� k                        8                                                                       ;�                      D                                                                      |��                     �                        �                                              }�                     ��                      �                                             }�?�                    ��                     �>                                             ;���                    D >                     ���                                            ���                   8 �                    ��                                            ^����                                         ^����                                          n���                    �                   .��                                           / ?���                                        / ?��                                          7���~                     �                  ���p                                          � ���                     p                  � ��                                          � ���                                       � ���                                         �  �>                     �                 �  �8                                         �  ���                     8                 �  ��                                         �   ��                                      �   ��                                        �   �<                     �                �   �0                                        �   �π                     0                �   ��                                        x    ?��                �                     x    ?�                                       x    �x                �     �               x    �`                                       �    ��                @      `                �    ��                                       �     ?�               @                      �     ?�                                        �     ��                                      ^     ��                                       �     �x                      �               ^     �`                                       o      �                      `               /      �                                       o      �                                    /      �                                       7�     ��                                    �     ��                                      7�     �x                     �              �     �`                                      �      �                      `              �      �                                      �      �                                   �      �                                      �      ��                                   �      ��                                     �      �x                     �             �      �`                                     �       �                      `             �       �                                     �       �                                  �       �                                     x       ��             �                     x       ��                                    x       �x             �        �            x       �`                                    �        �             @         `             �        �                                    �        �            @                      �        �                                     �        ��                                   ^        ��                                    �        �x                      �            ^        �`                                    o         �                      `            /         �                                    o         �                                 /         �                                    7�        ��                                 �        ��                                   7�        �x                     �           �        �`                                   �         �                      `           �         �                                   �         �  �                     �       �         �   p                               �         ��  p                  ��p       �         �� �                       `       �         �_���                  � �       �         �@ �                       �       �          ����                   @        �          � �                              �          ����                            �          � �                              x          ����        �                    x          � �                               x           ����        �             �       x           � t                               �           ?��r        @              r�       �           ���                               �           7� ��       @             ��       �           � w                               �           7� v                      7        ^           �                                �           7� 9�                     ?�       ^           � p                       0        o           7� A�                    ߠ       /           �  @                               o           7� `                    `       /           � 	�                      @       7�          7� �                    �       �          �                                7�          7� `                    �       �          �                                �          7� `                    7�       �          �                                 �          7� �                    �       �          � p                             �          7� `                    p       �          � �                              �          7� �                    �       �          �                                �          7�                     �       �          �                                 �          7�  �                    �       �          �  �                       �       x          7� �        �             �       x          �  `                       @       x          7�  �        �             �       x          � �                       �       �          7�         @            ~�       �          �                                 �          7�  9�       @             y�       �          �  '                       !        �          7�  t                      7�       ^          �                                 �          7�  0                      ?        ^          �  p                       0        o          7�   �                    ��       /          �  @                                o          7�  �                    o�       /          �                                 7�         7�  @                    �       �         �                                 7�         7�  @                    �       �         �                                 �         7�  �                    �       �         �                                 �         7�  �                    �       �         �                                 �         7�  �                    �       �         �  �                      �       �         7�  �                    �       �         �  �                       �       �         7�  �                    �       �         �   �                       �       �         7�                      D       �         �   �                       D       x         7�   �        �            �       x         �   �                       �       x         7�   Հ       �             �      x         �   �                       �       �         7�   ŀ��     @             �        �         �   � ��                    �       �         7�   ����     @             @        �         �                         @        �         7�   G���                          ^         �   8 >                             �         7�  ���                   �      ^         �    >                             o         ?� ����                  �       /          �   �>                             o         ?������                 �         /             ��                              7�        �������               �          �           �����                             7�        �����                �           �         ���                               �        �����                  .�            �        ���                                 �        ����                   .�            �        ��                                 �       ���                    .�            �       �                                   �       ��                                  �                                           ?����������             ��  �              8        �                                     �       ��             ?������              @�  � �                                      ����������               �  �                 ����������               �  �                 �������                                      ���������                                      ��������                                       ��������                                        �  �                  �  �                                                                 �                                              �                                              �    0                 �����                 �                                             ������                                        ������                                         �    <                                        �    4                                                                                                                                