�5l  Ȍ��                        x       �                                                  x       �                                                  x       �                                                  x       �                                                  � �    �                                                  � �    �                                                  � �    �                                                  � �    �                                                  � �    �                                                  � �    �                                                  � �    �                                                  � �    �                                                  ��<y��6�<�v���<                                              ��<y��6�<�v���<                                              ��<y��6�<�v���<                                              ��<y��6�<�v���<                                              y�f̀6ݳf�f���f                                              y�f̀6ݳf�f���f                                              y�f̀6ݳf�f���f                                              y�f̀6ݳf�f���f                                              �~���?ٿ~�f��~                                              �~���?ٿ~�f��~                                              �~���?ٿ~�f��~                                              �~���?ٿ~�f��~                                                                                                                                                                            �`���?ٰ`�f���`                                                                                                                                                                                                                                           ͛f́���f�f��sf                                                                                                                                                                                                                                           x�<x����<�f��c<�                                                                                                                                                                                                                                                         `                                                                                                                                                                                                                                                          �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ��          ��          ��          ��          ��                                                                                                                                                                                                      �"|         "'�        �"|         "'�        �"|          ݀          ��          ݀          ��          ݀          "           "           "           "           "                                                                         /���       ���<        /���       ���<        /���        � \          �        � \          �        � \                                                                                                                                   c�"~0       ?"'�        c�"~0       ?"'�        c�"~0        ݁�       ���        ݁�       ���        ݁�        "          "          "          "          "                                                                       �/���       ;���>�      �/���       ;���>�      �/���        A� \        �        A� \        �        A� \                                                                                                                             s���s�      �?���8      s���s�      �?���8      s���s�      �  �       �  �      �  �       �  �      �  �                                                                                                                         3�����`     9�����      3�����`     9�����      3�����`      `   1�      �         `   1�      �         `   1�          @                     @                     @                                                                      �����     �����{      �����     �����{      �����       �   @          �       �   @          �       �   @                    B                    B                                                                               �������     6������`    �������     �������    �������      f    0     	     �     f    0     `    3      f    0                  �    @                                                                                                         o�����v     M�������    o�����v     6������`    o�����v      �     �     2     `     �     �     	     �     �     �          D                      D     �    @         D                                                                    �������    ��������    �������     M�������    �������           &     D               &     2     `          &                        �                                                                                                         ��������   ��� ���    ��������   ��������    ��������    @           ��  @    @          D         @           �          �           �                �     �                                                                         >��� ����   �����    >��� ����   �������    >��� ����      �        �� $      �         �  @      �              �       �              �    �                 �                                                                   m��8 ����   ��  _���   m��8 ����   �����    m��8 ����      � � @   � p  ` 
      � � @     �� $      � � @       �        @ ���        �           �          �                                                                       ������X   ��� ����   ������X   ���_���   ������X    ( �  �    � �     ( �  �   � p�` 
    ( �  �      � �       1��`       � �      @ ��       � �                                                                    ���x ���   7��?����`  ���|���   ��ǀ���  ���x ���     ��� @    ?��  �    ��� @    ���      ��� @    @ �       �>�     @ �        8  �     @ �                                                                     ��� /��   k���) ����  ��� /��   7��8  ���`  ��� /��    � c� �0     �) ��@   � c� �0     ?��  �   � c� �0         �        �          �      �           �                                                                   ���  ���   w��� �p  ���  ��   k���  ���  ���  p��   @�� �     w� ` �  @��      �  �@  @�� �       `   0        � �       |   �         �        p  �                                                                  �    %��   ��� ����  �   E��   w��   _�p  �0 ���    �,  �    @ O ��    �  F     3� 8 ` �   �< �      �        0 � ` �    �   �        ��      � ��                     �            @                     �      ���   ��� o�� � ���  ��   ����  ���  `���  ��  �	���   �   y    �� �� H      �    @ C  ��    0 �	     � 0``      @ �      ��   �     <  ` �   �� ��                     �            �          `           �      ��    ��@ _�` � u��  ���   ���@ o��  � ���  ��   ��@  	 �   ��  �p � v (  	 �   ��  �� ��� H  	 ` 8���     0``      � �      �  �       x  � 0      � �                      �         �   �          �                  5��    �` ��� � ;��  5���  ��` _�H  '��  5�Ԁ ��`  
 7    @�  � � :   
 1�  �@�  �L  � (  
 4� >�@�   00`� � @  @  �     �  �� @   � �        � @                   �        �  �                            /��     ��� ��� � �  /���  ���� ���   ��  /�� � ?��   j    � @ @� � �   j�  �� @  �  2    i��   @   0`�`@      �      �  �@   @p �      �  �                    �         �  �                   �       [�     O�� �  � ��  [�v  ���� ��   ��  [� ?�� ���  $ �    �  �  � �
  $ �v  ��  @	      $ � ?�� �     `(a@�0       �       `�  �0     � �       n ?�� p                     �         v  �                   ?��      ���     /�X ��  � _�� ���;  po�X �    ��� ����}� O�X  (�     h �     � `  (�;� p� � �    �
  (��}� H �  @ @(aA@      �  �   @ @  �    � �     @ N��� 0                     �         ;  p                  �}�      ��@     �� 
��  � ��� ��@=  `7�� ��  @ �� ��V��� '��  @`     4 @  l  � �   @`=  `t @  7  @ @  @v��� $ @   �(����      �  @   �?� �   � � �   ����                     �         =  `                  ���     o��     �� �� �� ���o��� ��� ��  @ ?��o��������  ��        
 \ �� �   ��� �6   	 -  @     ������     
��� @      �        ?� � @   � �  �   ���� @                  �         � �                 ����    _�      �� �0 ��  ���_��� ��� ��      ��_������  �@        
 � ��  �   ��� �   
 R   @    �.���     
��     @  �  0     � �     !� �  �    ?����                    �         � �                  ���    ��  � 	� ?�� ��  k���� ���	� =�� �  ������?���   	� � 	�   � ��  l @  	��݀	�  � �\  � @  	.�?���   �

    @ �      � �    a� �  p   ��?�                    �         � �                  �>?�    ��  (� �� /�` ��  g���� h���� /�� �  _����<�����    *� � ` ��  d   j��� � �j  X  >����  @��4    � �     @ �߀    A�Ϝ  0   @�����         �        �         H ��        �       ���   ��  =�� �� +��  �  '���� }�� �� +�@ ��  '����<����� @  ?�� �  � ��  &  @ �� �  b ��  $  @>����@    ���H�     �       �߀�    ���      �����       �  �       �         \�  �      �        ���    �   � _� W��    2��� � � _� W�@  �  !���?� ��� �&  +�� `  (� ��  3  �& ��� `  (b ��  "  �&?����     B\Ȑ�             �� �   ���      ?�����        �  @                � �  @       �        ?� ��    �      � w�� e3  ��� � 6 � w��      ���?� ?��  �,  �� ` � ��     �, ��� ` � ��     �,?����`   �@  �     `2      � ?  �   �        ?�� ?� �            @               � 6  @                ?� ?� @  ��  &S  /����  g3  �x�� �S. /���� e2  �x���S?�/�� T  9�� 0 @� ��   � \ ��� 0 @ ��   � P����0  �!�R&4@h�    `2     �  �>  �   �`2     � ?��?� �        P                   �P.                �P?�    
��  fs0  �����     	�
��  �s<  ����� g3  ��
��??�s?� ��� X  y��  �  P� ��  	�  X  ��� �  P����   X??����@�     �I&(��`      �       �,  `    �`2       ��/��`        p                     �p,                ?�p/�    
��  ` 0  �����  �� ��
��  ` 0  �����  ���
���` 7� ��� X  ��  �  P  ��� �  X  ��  �  P���{�   X?�����     h%� �`      �        �   `    � ��     �� ��`       @           �         @           �     �@ �    �  ��<  W����  > � ���0 ��<  W����  ���� ���?��W��  � ���  X    >��� �P  � ���  �    ���E�P  �/������X  @� >� 0  P  ? �    @ � <  0  P � ���   @�� ?��0      � <        > �        � <         �     �� ?��  �� � >  _��_�  ?��� ?��� � >  _��_� > � E����/�� ?��_��
 � ���  X  �  ? � @ 
 � ���  �  � �>��� e� 
 �/������X    @	��  0     ~��� �   @ � ~  0    x? ���    @�� ��0      � >        > �        � >       > � A     �� ?��  �  ���  K��_�  ~� ?��  ���  K��_� ?��� ��� ?����o�K��
 0 � ~  L  �  �� @ 
 0 � ~  L  � ? � � 
 0?�� ~o�L    �O��� 8     ��y� �   � ���  8    ������   �������8      � >        | �        � >       > �  �    �� >o�  �@ �p? ���_�  ��� ��` �p?  +��_�  ~�<���@7��p??�+��
` �� �  �  � � @ 
` ��  l  � @��<
� 
`7���?��    �?�w��      ���� �   � �w��     ?��y���   ���w���      �         �  �        �         | �  �    �� ?�  �@ ������A��  ��� ���@ ��� /�A��  �������@{�����/�@ ` � ?����   ��� �( ` � ?� l�   � ���( `{�� ?��l�
 ���ό   � ��~| � 
 � ��π   � ���� �� 
 ��������      � �       �  x  �     � �       �  �  �    � ��  �@ �x�</��_� ��� ��@ �x� /��_� ��� B���@}πx��/��
` ���<,  � ꅊ�   
` ��� ,  � 0������ 
`}�����,    ���?w��     �z�| �   � ?w��     ��~| =�   ��?w����        �      � �<          �       �  x  �    �  ��  +�@ �8K��/��� ��B _�+�@ �8K� /��� 	��� ��+�@~^�8K߀/��` �X���, @ O�B ` ` �X�� , @ ꅊ� "� `~^�X���,    �x?W�W�     뿮�  �   � W�W�     �z�| �   ��W�W���       �        �   @      �      � �<  �     ^ ߀  +�� !8��< ���  �@ �+�@ !8��  ��� ��B _�+����8��>p�� � !D�<  @,  `@ `  @ !D�  6 @ O�B `  ���D�>q    瞻���     ��߾  �  � ����     뿮� �    ^���߈�        �          @   @       �          �   @     @ �    ?�� }�  ����  #�  �?�@ }�  ����  �@ _�?����}���� �   @ ,  4`` ` @   &@ ,  `@ 	` ����@ ~����  @ ˿�  � � >����  @ ��߾ �   >����l                      @                @   @          +�� >q�  ���  !ώ  _�+�  >q�  ���  #�  �+����>q��W��� F   @,  "�
  @   F   @,  4`` ` ���F�V    <����     ���  �  � <���� <    ˿� �    <����,                  G    @                      @           +�� ������  �_�( _�+�����������  !ώ  �+���������� ,p�� @,   H�  @ ���,p��� @,  "�
  ` ���,p��V    ���]�     ����  �  �����]���    ��� �    =��]�,       p          H�   @   ���p ��       G    @      p     +�� 
���?��� `_�4 _�+������������  �_�( �+��������7��� �� ? @,   H�  @ ������� @,   H�  ` ������v     =��}�     ����  �  �����}���    ����  �    =��}�       �          H�   @   ���� ��       H�   @      �     ?�� ��_������  �_�( _�?�  ��@ ���� `_�4 �?������G�7�� � ����@ ,   H�  @   ��  @ .   H�  ` ������6@?����}�  @ ����  � �����}��� @ ����  �   =��}�        �          H�   @      �          H�   @      �     +�� 
��� ���  !O�  _�+�  J��� ���  �_�( o�+����������� ��   @,  "�
  @   B��  @.   H�  p ������7   ? =��}�     ���  �  �����}���    ����  �    =��}�        �          G    @      �          H�   @      �     +�� �� ���  #�  �+�  B�� ���  !O�  o�+���������� ,p�  @,  $`  `   B,p�  @,  "�
  p ���,p��    �=��]�     ۿ��  �  �����]���    ���  �    =��]�        p               @      p          G    @      p     +�� :q� ���  �?@ �+�  :q�  ���  #�  o�+����:q����� F  @,  0 @ `   F  G @-  $`  p ���F�    �����     ��߾  �  � =���� <    ۿ��  �    =����                       @                      @            ?�� ������ �OB _�?�  �  ����  �?@ �?������� � �@ , PQB ` @   &@ .� 0 @ ` ����@  ~����  @ 믮�  � � >����  @ ��߾  �  ~����                        @                     @            +�� !=�<p��� �χ� ��+�  !=�  ��� �OB �+���=�/���� !E<p @ �ϋ� � @ !E   @/@PQB ` ���E?�    �����     �pu| �  � ����    �믮�  �   ^����                  �@<  �                       @             +�@ ��{��)��� � � ��+�@ ��{� )�����χ� ��+�X��{��)��` �����* @ ��� � @ ���� * @��ϋ� � z>�����*    �xWW�     ��~ �   � WW�    @�pu| �   � �WW�        �      �  8  �      �      �@<  �      �   �@ �p�?+��_� _���@���@ �p� +��_�� � �����^|o�p��+��
` ���?(  � _� �@� 
` ��� (  ������� 
|o����(    ���w��     ?������   � w��     ��}��   ��w��         �      �  �  �       �       �  8� �     �   �@ �����A��}~������@ ��� /�A��� �������O������/�@ ` � ��� }~����( ` � � ,� �� ���( ��� ��,�
 �����   � ���}��� 
 � ���   �����@� 
 �����       � �      || �� �     � �       �  �@ �   �� �   �@ �x?D /��_����������@ �x?  /��_�x~������G���x?y�/��
` ��?D ,  �������� 
` ��?  ,  ���~���� 
o����?y�,    � o�w߀    �~z����   � �w߀    8��}� �   �~�w߆       �       �> ��� �     �        | �  �     �     �  �8�� K��_���`7�=���  �8�  K��_�>��������#���8�|�K��
0 �X�� L  �	��`7��� 
0 �X�  L  �~������ 
7���X���L    � ��?  8   �?���~    � �?  8   �~z���   � �? 8      �>      � �<      �>        > ��  �     �>    �� �~I�W��_�_O����}���� �~  W��_���`7��������~�`W��
 � �~I�P  �_�����}� 
 � �~  P  �?��`7��  
 �����`P    @���  8   ���?��    @ ���  8     ?����   @ ����8      � ~       ��      � ~         �       � ~    �� s���&@_����}>������� ���  _������������������� _��  � s���&@X  }������P  � ���  X  �������P  ������� X  @��  0  P� ����   @ ��  0  P  �?�   @ �� �0      ��      | �� �      ��        ��       ��    
�P���!������t��� ����
�P  ��  �������� �
�
�P������ ����!��  Pw�����   �  ��  �  P�����
�  �?������     0 ���  p   � �� �       ���  p     ���      ��� @p       ��       p ��  �       ��         ��         ��     
�P	���P������� �� >3��
�P ?��  �����  �� |��
�P ������� �	���P�  P�� �� �   � ?��  �  P���� �   ��������     � ?��  `     ��  ~       ���  `     ��        ?��  `       ?��          ��  2       ?��         ��         ?��     ���O��H9/����� _� ��x��  /�� /�����  �� <�x�� ?�����/�� \�O��H90 @�� ]� � � \  /�� 0 @� �� } � \?ﯟ��0  �!  ��  �     ?�  >   �  ���  �    ��    �  ���  �       ��          �         /��          ��         ��     � $M�R$_� w��     ����  E�	 _� w��  _� <������?��_�  �o $M�R$@ �     �   �l  E�	 @ �  �� =   �l���?��@    �   �          <    ��~  �      ?�      �   �       �   @                  A�  @       �         �   @  � X��I� W�|     ���� � D � W��  � '�����<���� �. X��I`  (|     �  �. � D `  (�  #� =&  �.��>���`          �    �      8     � ? �              �  !�            @                  �   @                       @  �� ��)
�� +��     �����  � ��� +�`  � )����������� @6 ��)
�  �     �  @6  � ��  `  � ?*  @6������          �    @      8     � ? �    �               �            �                  �   �                       �  ��A$�%� -��     ����� 	  " � /�0  � W���� �������  A$�%@  �     �   	  " @ 0  � T   ������@  @      �   @      p   @ � ��   �     8   @      �                       0                                   ����E(����� =��     ?�����  @	�� =��  � ������������   	��E(����  l     0 @  	�  @	�  �  � � @  	�������            0      �    � �    `     p                                                                     _���(���� ��     O��_��   � �L  � ���_��������  ���(����  	 t     P   ��   �  
 �  � �   ��?������                     �     � �     0     p                                @                                    o�l
(����� ��     ���o�`$   �5�� ��  � _��o�`�������  �l
(���    
     �  �`$   �5   	 v  � ?P   �`�����     �               �    �� �          �    �                          �        �           @              ���

(�@k�� ��     ?�� ����  �k�� ��  � ��� ���������  @�

(�@j @       @   @��  �j @  +  � >�  @����� @   �               �    �?  �         �    �          �                     �   �           �     �         ��P(`���� ���    ��� ��PH  @��� ��    =�� ��P������   P(`��    �        XH  @�      /� =@   P����     �     8                �?  �8         �     �    8      @                     @   @                @         �,(`���� ��@    $��  �,�   )��� ���   z��  �, ;�����    �(`��    @`    %     ��   )�     
� _  z�     � ;���      p     p     �          p~  �p                p    p                                                              ;��(`c_�� ���    K��  ;��  #_�� ��` >  u��  ;�� � _��   V(`cP    �    H    W  #P   @` �  �    V � P     8     �     �    <      8�  ��     � @        8    �           @      �              @                     @    /��00P$��` ��L   ���  /��"   ��` ��� |  ���  /�� � ��`   )00P$� �   L   �     ("   � �  �| �    )�� � �        �      �    x      �  ��     � �  <         �           �      @              �      �               �    ���009��  ���   o�x  ��   �� ��L � ���  ���� ��    �009@     s   ` �       @     M�� �      �π 9@          �      <   �      �   ��      �   x       0  �                 0    `                 @                   �000f���  _���  ���  �  ���  ����� o�x  �>?  f���   �000f�     (�  �     �  �    3�� h �   �>?  f�     �             �      �   �       |�  �      ��                        �                 0�   `              ���001���   ��8  ����  ���  	��   _���� ���  ���� ���    �001�      8  �     �  	      )�� �     �� �      �   >       �         �   �          �      �   >        �                     �              �       �        ��c�0>=��   =��ǀ���  ��a� =��   ��?  ����  ��c� =��      c�0>>      ǀ       a� >>       ?� ��       c� >        �  �       �  �        �  �       �          �  �        `   0       �          `   0                  `   0     ���x0����   ����{���  ���x ����   =��ǀ��  ���x ����      x0��      ��|       ~��      ǀ�      x ��        ?� �        ��        ?� �       �  �        ?� �          �        0  `          �       �            �     �������   ��߀���  �������   ����k���  �������    @ ��     @ ?��     @ ��      ��l     @ ��       � �         ���        � �         ��        � �                    ��                   0  `                 ���� ����   ��������    ���� ����   ������   ���� ����     � �        ��        � �      @ /��      � �        ���          �         ���         ���        ���          � �          �          � �         ��         � �       ����o���   �������    ����o���   �������    ����o���       g�p       �  �         g�p         �          g�p          ��                      ��         ��          ��          �                       �           �          �        7�������`   �������|    7�������`   �������    7�������`      �   �          �      �   �    �  �        �   �                                                                                                                                  �������    �������    �������   �������|    �������     �                       �                �     �                                                                                                                                        �������     .�������    �������     �������    �������                       @                                                                                                                                                                        ������z     �������    ������z     .�������    ������z          �                      �          @         �                                                                                                                                   �������     ������     �������     �������    �������                      D                                                                                                                                                                          ^������     ������      ^������     ������      ^������      !    @         D      !    @         D      !    @                                                                                                                                    ?������     ������      ?������     ������      ?������          @                     @                     @                                                                                                                                     ������      ������      ������      ������      ������                                                                                                                                                                                       �����       =�����      �����       =�����      �����                                                                                                                                                                                             }����       ����        }����       ����        }����        "          "          "          "          "                                                                                                                                       ����       ����        ����       ����        ����                                                                                                                                                                                                 ���         ���        ���         ���        ���          "           "           "           "           "                                                                                                                                         ��          ��          ��          ��          ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               �         �          ` �       �          `  `                                                                                                                                                                                                    0         �  <        ` 0       �  3        `  �                                                                                                                                                                                                              �          �  0       �          �  �                                                                                                                                                                                                    Ǜ>       �x�        珀0       �x�        珁�                                                                                                                                                                                                    �l�3f       ��        �ـ`       ��        �ف�                                                                                                                                                                                                     6l�?f       �}�        �ـ�       �}�        �ك`                                                                                                                                                                                                     6l�0f       �͘        lف�       �͘        lك�                                                                                                                                                                                                    6l�3f       �͘        lك        �͘3        lـ`                                                                                                                                                                                                    �Ǚ�>       �|�        gσ�       �|�        gπ`                                                                                                                                                                                                                              �                      �                                                                                                                                                                                                                   �                      �                                                                                