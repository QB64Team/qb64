�d  �~                       �      �    0    �                                              �      �    0    �                                              �      �    0    �                                              �      �    0    �                                             3 � `    �       �                                             3 � `    �       �                                             3 � `    �       �                                             3 � `    �       �                                             0 � `    �       �                                             0 � `    �       �                                             0 � `    �       �                                             0 � `    �       �                                             0<�p<�6��3�7ǀ�6�                                             0<�p<�6��3�7ǀ�6�                                             0<�p<�6��3�7ǀ�6�                                             0<�p<�6��3�7ǀ�6�                                             fٳ`���6��l��6ـ                                            fٳ`���6��l��6ـ                                            fٳ`���6��l��6ـ                                            fٳ`���6��l��6ـ                                            ~߰`>����3�o��6߀                                            ~߰`>����3�o��6߀                                            ~߰`>����3�o��6߀                                            ~߰`>����3�o��6߀                                                                                                                                                                              `�0`f�͛1��l f6�                                                                                                                                                                                                                                                3fٳ`f��͛v��l��ـ                                                                                                                                                                                                                                               <�0>�6���7ǀ��6�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               p                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       �                                           �                  �                                           �                  �                                           �                  �                                           �                                                                                   �                                            �                   �                                           �                                                                                  ?�                                          ?�                 ?�                                          ?�                  ��                                           ��                  ?�                                           ?�                  ��                                           ��                 ��                                          ��                 ��                                          ��                  ��                                           ��                 ��                                          ��                 ��                                          ��                 ��                                          ��                 ��                                          ��                                                                              �                                          �                 �                                           �                                                                                                                                                .`                                           .`                  ��                                          ��                                                                                !�                                          !�                 ]��                                          ]��                 >@                                           >@                                                                                 Z�                                           Z�                  Z�                                           Z�                  =                                            =                                                                                  1                                            1                   ��                                           ��                  |                                            |                   0                                            0                   2                                            2                   �                                            �                   x                                            x                   0                                            0                   �                                            �                   �                                            �                   x                                            x                   `                                            `                   l                                            l                   n                                            n                   �                                            �                   `                                            `                   d                                            d                   n                                            n                   �                                            �                   `                                            `                   d                                       �   d                   l                                       �   l                   �                                            �                   `                                            `                   d                                         d                   l                                      ~   l                   �                                      �   �                   `                                           `                   ,                                     ��   ,                   ,                                     ��   ,                   �                     �                �   �                                                           �                       �                     �               |�   �                   �                     3�              ��   �                   p                     �               ��   p                                         �                �                       �                     �              ��   �                   �                     O�              ��   �                   p                     ?�               ��   p                                         �               �                       ,                     <              ��   ,                   �                     �             ��   �                   p                     �              ���   p                                         <               �                       |                     q              �    |                   �                    q�             ?�    �                   0                     �               ����   0                   0                     p               �     0                   R                     �             ����   R                   V                    �             ����   V                   8                    ��             ���    8                                        �               ��                        R                    �            � p   R                   V                    ۘ            >� �   V                   8                    �             ����    8                                       �              �                                             �            ��                         W                    �            �� ��   W                   8                    �             ���     8                                       �             �                          >                                ���   >                                       8   ����    |����                                          �            ���                                                           �                          )                        ����   �� x�    )                   +                    p   ����   �� ���   +                                       �            ?���                                                          �                           )                    @           x?� �     )                   +                    `          �?����    +                                       �   �8�   ���                                                           ?�                                               �          ���?                         +�                   �          ?�����     +�                                          A   ��                                                           �                                                @  �A   �p�                         ?�                   � �A  ���      ?�                                         �����������                                                   A   �                            �                   @ �����������       �                  �                   � ������������       �                                        �����������                                                   ����������                             �                   @ ����������        �                  �                   � �����������        �                                        ��y�y����                                                   ��y�y���                              �                   �  ��~  =��         �                  �                   � / ��~  ?���        �                                        ��8����                                                                                           �                     @��>  ~          �                  �                   � \����������         �                                      @ ?�                                                                                                   �                   � 8���>  ~           �                @�                   � ����>  �          �                �                    @ ~�}�����                                                   8                                       
@                     t��}��              
@                �
�                    v�                   
�               �                    � ����>                               @                       p                                       
@                     j  <��              
@               `
�                   k  @              
�               `                    � � ��~                               ��                       `  @                               @@                   � ����              @              ��`
�                   
� ����              
�              ��`                    ��                                    ��                       �                                     �@�                   �� ����              �              <� �                   ��                    �              ��`                    p� ����                             ���                      �                                    �                      �`                                  ��  p                   �;t                    p             �� `�                   <�                    �              ?���                                                         �  `                    f�                    `             x?� �p                   ��                    p            �?� ��                   �                    �             ���                                                          ?�  �                    1�                    �            ��  �                   q��                    �            �� ��                    ��                     �             ���  �                    �                      �             �   x                                         x            ��� |                    ��                    |           �����                    C�@                    �            ���   @                                            @             �   <                    #��                    <           � p  >                    o��                    >           ?� �� �                                          �            ����                                                             �    �                                         �           ��� ��                    3��                    �          ������ p                                          p           ���                                                            ��     �                                          �          ��� ��                                        ��         ~����                      �                                ���                                                            �      w�        �����                             w�        �� p�   ��        �����                             ��        �� ��                                                         ?���                                                           �       -�                                           -�        ?��    }��                                          }��      �?���    �        �����                             �        ���      �                                           �         ?�       �����������������                          �����������     ?�����������������                          ?��������#����     �        �����                              �       ���        p        �����                              p        �        ��       �����                             ��      ��@?      ��       �����                             ��      ����      ?�����������������                           ?�����������        �       �����                              �      ��        ?����������������                          ?���������      �?����������������                          �?����������       �����������������                           ����������          ?����������������                            ?��������          ��                                           ��      ��       ��                                          ��      ���         ?����������������                            ?�������                                                                            �                                           �       �         ���������    ���                           ����������                  �����                                                                                                                    ����������������                            ��������          �����������������                           ����������                                                                                                                                                                                                                     �����                                                                                                                                                                                             �����                                                           �����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �0   3`        1�  ��    �          0                                                                                                                                                                                                                       `  0`  f`        1�  �    �          0    f                                                                                                                                                                                                                    `  0`  f`        1�  �    �          0    f                                                                                                                                                                                                                6�w<Ͼp3wg�       1���?�<���ǀ       0<��w��<|��ǟ                                                                                                                                                                                                        ��fٻ`m�fl�       ?�n����6ٳ��7l�       0f��g`�f�7lݳ                                                                                                                                                                                                        ��f>ٳ`m�fo�       1�l��٘6߳>͛6o�       0f��f`�~��6lٿ                                                                                                                                                                                                        ��ffٳ`m�fl       1�l��٘6�3f͛6l        0f��f`�`͛6lٰ                                                                                                                                                                                                        ��ffٳ`m�fl�       1�l��٘6ٳf͛6l�       0ff3f`�f͛6lٳ                                                                                                                                                                                                        ��6>ϳ0m�fg�       1����͘6�>���g�       ?<f36`�<|��g��                                                                                                                                                                                                              �               `       �                                                                                                                                                                                                                                                      �      > �                    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      A      P                                                                                                                                                                                                                                                           A  @   H                                                                                                                                                                                                                                                           A  @   H                                                                                                                                                                                                                                                         9c�c�`z'3�                                                                                                                                                                                                                                                         �A�A@� �H                                                                                                                                                                                                                                                         =A�@�'�H                                                                                                                                                                                                                                                         EA@�(�H                                                                                                                                                                                                                                                         EAQ@�h�H                                                                                                                                                                                                                                                         =�� y���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �                                                                                               