��e  ') . ������      ������      ������  �  ������  �  ������  ?�  ������  ?�  ������  ��  ������  ��  ������ ��  ������ ��  ������ ��  ������ ��  ������ ��  ������ ��  ������ ?��  ������ ?��  ������ ?��  ������ ?��  ������ ?�  ������ ?�  ������ <�  ������ <�  ������ 0�  ������ 0�  ������  �  ������  �  ������  �  ������  �  ������  �  ������  �  ������  �  ������  �  ������  �  ������  �  ������  �  ������  �  ������  �  ������  �  ������      ������  �  ������      ������  �  ������      ������  �  ������      ������  �  ������      ������  �  ������      ������  �  ������      ������  �  ������      ������  �  ������      ������  �  ������      ������  �  ������      ������  �  ������      ������  �  ������      ������  �  ������      ������  �  ������      ������  �  ������      ������      ������      ������      ������      ������      ������      ���������p ������      ������� � ������      ������D  ������      ������D  ������      �������'� ������      ������$   ������      ������� @ ������      ������ � ������      ������ �   ) . ������ ��  ������ ��  ������ ��  ������ ��  ������ ?��  ������ ?��  ������ ��  ������ ��  ������ ���  ������ ���  ������ �   ������ �   ������� ?  ������� ?  ������� ?� ������� ?� ������� � ������� � ������� � ������� � ������� � ������� � ������   � ������   � ������   � ������   � ������   ?  ������   ?  ������     ������     ������   ~  ������   ~  ������   �  ������   �  ������  �  ������  �  ������  �  ������  �  ������      ������  �  ������      ������  �  ������      ������  ?�  ������      ������  �   ������      ������ �   ������      ������ �   ������      ������ �   ������      ������ ?�   ������      ������ ��   ������      �������    ������      �������    ������      ���������� ������      ���������� ������      ���������� ������      ���������� ������      ������      ������      ������      ������      ������      ������      �������� ������      ������B�  ������      ������E�  ������      ������E�  ������      �������� � ������      ��������  ������      ��������  ������      ������P�  ������      ������P��   ) . ������ ��  ������ ��  ������ ��  ������ ��  ������ ��  ������ ��  ������ ���  ������ ���  ��������  ��������  �������   �������   ������� ?� ������� ?� ������� � ������� � ������� � ������� � ������   � ������   � ������   � ������   � ������   � ������   � ������   ?  ������   ?  ������     ������     ������  �  ������  �  ������  ��  ������  ��  ������  ��  ������  ��  ������  ��  ������  ��  ������  ��  ������  ��  ������      ������   �  ������      ������   ?� ������      ������   � ������      ������   � ������      ������   � ������      ������   � ������      ������� � ������      ������� � ������      ������� � ������      ������� � ������      ��������  ������      ���������  ������      ������ ���  ������      ������ ?��  ������      ������ ��  ������      ������      ������      ������      ������      ������      ������      ������� @ ������      ������B�� ������      ������E�� ������      ������E�@ ������      ��������@ ������      ��������@ ������      ��������� ������      ������P�@ ������      ������P�@   ) . ������      ������      ������  �  ������  �  ������  �  ������  �  ������  �  ������  �  ������  �  ������  �  ������  ?�  ������  ?�  ������  �  ������  �  ������  ��  ������  ��  ������ ��  ������ ��  ������ ��  ������ ��  ������ ��  ������ ��  ������ ��  ������ ��  ������ ��  ������ ��  ������ ?�  ������ ?�  ������ �  ������ �  ������ ��  ������ ��  ��������  ��������  ��������  ��������  ��������  ��������  ������      ��������  ������      ��������  ������      ��������  ������      ���������� ������      ���������� ������      ���������� ������      ���������� ������      ������  �  ������      ������  �  ������      ������  �  ������      ������  �  ������      ������  �  ������      ������  �  ������      ������  �  ������      ������  �  ������      ������      ������      ������      ������      ������      ������      ������� @ ������      ������B�� ������      ������E�� ������      ������E�@ ������      ��������@ ������      ��������@ ������      ��������� ������      ������P�@ ������      ������P�@   ) . ������      ������      ���������  ���������  ���������  ���������  ���������  ���������  ���������  ���������  �������    �������    �������    �������    �������    �������    �������    �������    �������    �������    �������    �������    ���������  ���������  ���������  ���������  ���������  ���������  ���������  ���������  ��������  ��������  ������� � ������� � ������� ?� ������� ?� ������� � ������� � ������      ������� � ������      ������   � ������      ������   � ������      ������   � ������      ������   � ������      ������   � ������      ������� � ������      ������� � ������      ������� ?� ������      �������   ������      ��������  ������      ���������  ������      ������ ���  ������      ������ ?��  ������      ������ �   ������      ������      ������      ������      ������      ������      ������      ������� @ ������      ������B�� ������      ������E�� ������      ������E�@ ������      ��������@ ������      ��������@ ������      ��������� ������      ������P�@ ������      ������P�@   ) . ������ ��  ������ ��  ������ ��  ������ ��  ������ ��  ������ ��  ������ ?��  ������ ?��  ������ ��  ������ ��  ������ � � ������ � � ������� � ������� � ������� � ������� � ������� � ������� � ������� � ������� � �������    �������    �������    �������    ��������  ��������  ���������  ���������  ���������  ���������  ���������  ���������  ���������� ���������� ������� ?� ������� ?� ������� � ������� � ������      ������� � ������      ������� � ������      ������� � ������      ������� � ������      ������� � ������      ������� � ������      ������� � ������      ������� � ������      ������� � ������      ������� ?� ������      ������ ���� ������      ������ ��  ������      ������ ?��  ������      ������ ��  ������      ������ ��  ������      ������      ������      ������      ������      ������      ������      ��������� ������      ������!A ������      ������"�@ ������      ������"�@ ������      �������O�  ������      ������H@@ ������      �������@� ������      ������(A  ������      ������(A�   ) . ������      ������      ���������� ���������� ���������� ���������� ���������� ���������� ���������� ���������� ������   � ������   � ������   � ������   � ������   � ������   � ������   ?  ������   ?  ������     ������     ������   ~  ������   ~  ������   �  ������   �  ������   �  ������   �  ������  �  ������  �  ������  �  ������  �  ������  �  ������  �  ������  �  ������  �  ������  �  ������  �  ������  �  ������  �  ������      ������  �  ������      ������  �  ������      ������  �  ������      ������  ?�  ������      ������  ?   ������      ������     ������      ������  ~   ������      ������  �   ������      ������  �   ������      ������ �   ������      ������ �   ������      ������ �   ������      ������ �   ������      ������ �   ������      ������ �   ������      ������      ������      ������      ������      ������      ������      ��������� ������      ������!A ������      ������"�@ ������      ������"�@ ������      �������O�` ������      ������H@ ������      �������@ ������      ������(A ������      ������(@�   ) . ������ ��  ������ ��  ������ ��  ������ ��  ������ ��  ������ ��  ������ ���� ������ ���� ������� � ������� � ������� � ������� � ������� � ������� � ������� � ������� � ������� � ������� � ������� � ������� � ������� � ������� � ������� � ������� � ������� ?� ������� ?� ������ ���� ������ ���� ������ ?��  ������ ?��  ������ ��  ������ ��  ������ ��  ������ ��  ������ ��  ������ ��  ������ ���� ������ ���� ������      ������� � ������      ������� � ������      ������� � ������      ������� � ������      ������� � ������      ������� � ������      ������� � ������      ������� � ������      ������� � ������      ������� � ������      ������� � ������      ������ ���� ������      ������ ��  ������      ������ ��  ������      ������ ��  ������      ������      ������      ������      ������      ������      ������      ��������� ������      ������!A ������      ������"�@ ������      ������"�@ ������      �������O�` ������      ������H@ ������      �������@ ������      ������(A ������      ������(@�   ) . ������ ��  ������ ��  ������ ��  ������ ��  ������ ?��  ������ ?��  ������ ���  ������ ���  ��������  ��������  ������� � ������� � ������� ?� ������� ?� ������� � ������� � ������� � ������� � ������� � ������� � ������� � ������� � ������� � ������� � ������� � ������� � ������� � ������� � ������� � ������� � ������� ?� ������� ?� ������� � ������� � ���������� ���������� ������ ���� ������ ���� ������      ������ ��� ������      ������ ��� ������      ������ �� ������      ������   � ������      ������   � ������      ������� � ������      ������� � ������      ������� ?� ������      ������� ?� ������      ������� �  ������      ������ ���  ������      ������ ��  ������      ������ ?��  ������      ������ ��  ������      ������ ��  ������      ������      ������      ������      ������      ������      ������      ��������� ������      ������!A ������      ������"�@ ������      ������"�@ ������      �������O�` ������      ������H@ ������      �������@ ������      ������(A ������      ������(@�             