��Z  �^r� �����������������������������������������������                                               �����������������������������������������������������������������������������������������������                                             @                                               �                                             @�                                             @����������������������������������������������@                                               ����������������������������������������������@����������������������������������������������@�                                            @                                               �                                            @�                                            @�                                            @                                               �                                            @�                                            @�                                            @                                               �                                            @�                                            @�                                            @                                               �                                            @�                                            @�                                            @                                               �                                            @�                                            @�                                            @                                               �                                            @�                                            @���������������������������������������������@ �������������������������������������������� ���������������������������������������������@�                                            @�@                                           �@ @                                           � �@                                           �@�                                            @�@                                           �@ @                                           � �@                                           �@�                                            @�@                                           �@ @                                           � �@                                           �@�                                            @�@                                           �@ @                                           � �@                                           �@�                                            @�@                                           �@ @                                           � �@                                           �@�                                            @�@                                           �@ @                                           � �@                                           �@�                                            @�@                                           �@ @                                           � �@                                           �@�                                            @�@                                           �@ @                                           � �@                                           �@�                                            @�@                                           �@ @                                           � �@                                           �@�                                            @�@                                           �@ @                                           � �@                                           �@�                                            @�@                                           �@ @                                           � �@                                           �@�                                            @�@                                           �@ @                                           � �@                                           �@�                                            @�@                                           �@ @                                           � �@                                           �@�                                            @�@                                           �@ @                                           � �@                                           �@�                                            @�@                                           �@ @                                           � �@                                           �@�                                            @�@                                           �@ @                                           � �@                                           �@�                                            @�@                                           �@ @                                           � �@                                           �@�                                            @�@                                           �@ @                                           � �@                                           �@�                                            @�@                                           �@ @                                           � �@                                           �@�                                            @�@                                           �@ @                                           � �@                                           �@�                                            @�@                                           �@ @                                           � �@                                           �@�                                            @�@                                           �@ @                                           � �@                                           �@�                                            @�@                                           �@ @                                           � �@                                           �@�                                            @�@                                           �@ @                                           � �@                                           �@�                                            @�@                                           �@ @                                           � �@                                           �@�                                            @�@                    �               �      �@ @                    �               �      � �@                    �               �      �@�                                            @�@   > �@�    c c�  �      �`����   �@ @   > �@�    c c�  �      �`����   � �@   > �@�    c c�  �      �`����   �@�                                            @�@  � ���  ?� c g0  ?�      �`���   �@ @  � ���  ?� c g0  ?�      �`���   � �@  � ���  ?� c g0  ?�      �`���   �@�                                            @�@  � �À  p  � �0  |p        �0 >   �@ @  � �À  p  � �0  |p        �0 >   � �@  � �À  p  � �0  |p        �0 >   �@�                                            @�@   �� ��  �  � �`  0      ` �`    �@ @   �� ��  �  � �`  0      ` �`    � �@   �� ��  �  � �`  0      ` �`    �@�                                            @�@   �� ��  6�  ��`  0      `�0`    �@ @   �� ��  6�  ��`  0      `�0`    � �@   �� ��  6�  ��`  0      `�0`    �@�                                            @�@   �� �>  6  ���  0      ��0@ <   �@ @   �� �>  6  ���  0      ��0@ <   � �@   �� �>  6  ���  0      ��0@ <   �@�                                            @�@  � �|  f  3���  0fc�����0 ���   �@ @  � �|  f  3���  0fc�����0 ���   � �@  � �|  f  3���  0fc�����0 ���   �@�                                            @�@  > 1��  ��c�   '���?���0`��?�   �@ @  > 1��  ��c�   '���?���0`��?�   � �@  > 1��  ��c�   '���?���0`��?�   �@�                                            @�@  �0 ϐ ����1�   �����0a�0 &    �@ @  �0 ϐ ����1�   �����0a�0 &    � �@  �0 ϐ ����1�   �����0a�0 &    �@�                                            @�@  �0��0 ����0�   p30� ��  c    �@ @  �0��0 ����0�   p30� ��  c    � �@  �0��0 ����0�   p30� ��  c    �@�                                            @�@                                           �@ @                                           � �@   `��` f03 �   �&8�  � ` �    �@�                                            @�@                                           �@ @                                           � �@   `�` 0`�0� �|�<  � ` ��   �@�                                            @�@                                           �@ @                                           � �@   ��� 0`� � ��<��  � ���   �@�                                            @�@                                           �@ @                                           � �@   ��� 00�x   �0��g�   ��`   �@�                                            @�@                                           �@ @                                           � �@  ��� `8~0�x�  �0���  � 0   �@�                                            @�@                                           �@ @                                           � �@  �0�� ��`�0�   `��� ?�0��    �@�                                            @�@                                           �@ @                                           � �@  �`� ����1�   `���� ?�0��    �@�                                            @�@                                           �@ @                                           � �@                        ��             �@�                                            @�@                                           �@ @                                           � �@                                         �@�                                            @�@                                           �@ @                                           � �@             0                             �@�                                            @�@                                           �@ @                                           � �@             0                             �@�                                            @�@                                           �@ @                                           � �@             `                             �@�                                            @�@                                           �@ @                                           � �@                                           �@�                                            @�@                                           �@ @                                           � �@                                           �@�                                            @�@                                           �@ @                                           � �@                                           �@�                                            @�@                                           �@ @                                           � �@                                           �@�                                            @�@                                           �@ @                                           � �@                                           �@�                                            @�                                            @�                                            @ @                                           � �                                            @�                                            @�                                            @ @                                           � �                                            @�                                            @�                                            @ @                                           � �                                            @�                                            @�                                            @ @                                           � �                                            @�                                            @�                                            @ @                                           � �                                            @�            `�                              @�            `�                              @ @           `�                              � �                                            @�       >���  �          @0            @�       >���  �          @0            @ @      >���  �          @0            � �                                            @�       ���0  ?�          �0            @�       ���0  ?�          �0            @ @      ���0  ?�          �0            � �                                            @�      �0  |p          �`    0        @�      �0  |p          �`    0        @ @     �0  |p          �`    0        � �                                            @�      ��0`  0         �`     0        @�      ��0`  0         �`     0        @ @     ��0`  0         �`     0        � �                                            @�       �0`  0         ��              @�       �0`  0         ��              @ @      �0`  0         ��              � �                                            @�       �0 �  0         ��     `        @�       �0 �  0         ��     `        @ @      �0 �  0         ��     `        � �                                            @�       �0`�  0fc��� Bs�! @<      @�       �0`�  0fc��� Bs�! @<      @ @      �0`�  0fc��� Bs�! @<      � �                                            @�       � `   '���?� 8�0��c<| |��>      @�       � `   '���?� 8�0��c<| |��>      @ @      � `   '���?� 8�0��c<| |��>      � �                                            @�      �<`�   ���� ܶ1�<b�� �ǆf      @�      �<`�   ���� ܶ1�<b�� �ǆf      @ @     �<`�   ���� ܶ1�<b�� �ǆf      � �                                            @�      0�x`�   p30��a��Ǚ���<�      @�      0�x`�   p30��a��Ǚ���<�      @ @     0�x`�   p30��a��Ǚ���<�      � �                                            @�                                            @�                                            @ @     0����   �&8� 9�c�'��381� �      � �                                            @�                                            @�                                            @ @     0Ca���0� �|�< s�ǈ��60���      � �                                            @�                                            @�                                            @ @     0Fg0�  � ��<�� s��1�dp�;�      � �                                            @�                                            @�                                            @ @     0n�1�    �0��g� 1��3l�3?      � �                                            @�                                            @�                                            @ @     |�a� �  �0��� 3f1�c��bp:0      � �                                            @�                                            @�                                            @ @     9�c �   `��� >L3�8f0���`��      � �                                            @�                                            @�                                            @ @     ����   `���� �aF1�����      � �                                            @�                                            @�                                            @ @       @         ��         �  ?        � �                                            @�                                            @�                                            @ @                            !�           � �                                            @�                                            @�                                            @ @                        0    1�           � �                                            @�                                            @�                                            @ @                        0    3�           � �                                            @�                                            @�                                            @ @                        `    3            � �                                            @�                                            @�                                            @ @                         `                � �                                            @�                                            @�                                            @ @                         �                � �                                            @�                                            @�                                            @ @                         �                 � �                                            @�                                            @�                                            @ @                         �                 � �                                            @�                                            @�                                            @ @                                           � �                                            @�                                            @�                                            @ @                                           � �                                            @�                                            @�                                            @ @                                           � �                                            @�                                            @�                                            @ @                                           � �                                            @�                                            @�                                            @ @                                           � �                                            @�                                            @�                                            @ @                                           � �                                            @�                                            @�                                            @ @                                           � �                                            @�                                            @�                                            @ @                                           � �                                            @�                                            @�                                            @ @                                           � �                                            @�                                            @�                                            @ @                                           � �                                            @�                                            @�                                            @ @                                           � �                                            @�                                            @�                                            @ @                                           � �                                            @�                                            @�                                            @ @                                           � �                                            @�                                            @�                                            @ @                                           � �                                            @�                                            @�                                            @ @                                           � �                                            @�                                            @�                                            @ @                                           � �                                            @�                                            @�                                            @ @                                           � �                                            @�                                            @�                                            @ @                                           � �                                            @�                                            @�                                            @ @                                           � �                                            @�                                            @�                                            @ @                                           � �                                            @�                                            @�                                            @ @                                           � �                                            @�                                            @�                                            @ @                                           � �                                            @�                                            @�                                            @ @                                           � �                                            @�                                            @�                                            @ @                                           � �                                            @�                                            @�                                            @ �������������������������������������������� �                                            @�                                            @�                                            @                                               �                                            @�                                            @�                                            @                                               �                                            @�                                            @�                                            @                                               �                                            @�                                            @�                                            @                                               �                                            @�                                            @�                                            @                                               �                                            @�                                            @�                                            @                                               �                                            @����������������������������������������������@����������������������������������������������@                                               ����������������������������������������������@�                                             @�                                             @                                               �                                             @����������������������������������������������������������������������������������������������                                               �����������������������������������������������