�4a  XZA� �����������������������������������������                                                                                                                           �����������������������������������������                                                                                                                           �����������������������������������������                                                                                                                           �����������������������������������������                                                                                                                           �����������������������������������������                                                                                                                           �����������������������������������������                                                                                                                           �                                      ����������������������������������������                                                                                   ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀           � `       �                         � `       �                         � `       �             ���������������������������������������߀           �         �`                        �         �`                        �         �`            ���������������������������������������߀         �  �         �`                      �  �         �`                      �  �         �`            ���������������������������������������߀          ��7ͱ�g�Ͱ<y���s�                      ��7ͱ�g�Ͱ<y���s�                      ��7ͱ�g�Ͱ<y���s�           ���������������������������������������߀          a�6m�0m��m�fͶͳf`                      a�6m�0m��m�fͶͳf`                      a�6m�0m��m�fͶͳf`           ���������������������������������������߀          a�6m��f6o�`ͶͿg�                      a�6m��f6o�`ͶͿg�                      a�6m��f6o�`ͶͿg�           ���������������������������������������߀          a�6m� c6o�`ͶͰf                       a�6m� c6o�`ͶͰf                       a�6m� c6o�`ͶͰf            ���������������������������������������߀          a�vm�0m�6f`fͶͳf`                      a�vm�0m�6f`fͶͳf`                      a�vm�0m�6f`fͶͳf`           ���������������������������������������߀          `��͙�g3�`<y���3�                      `��͙�g3�`<y���3�                      `��͙�g3�`<y���3�           ���������������������������������������߀                         �                                        �                                        �              ���������������������������������������߀                         �                                        �                                        �              ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ������������������������������߿�����߀                                                                                   �          �     @A      @     ���w����������������������������������߀                                                                                    �     �           @A      @     ���w����������������������������������߀                                                                                    �     �           @A      @      ���t�1�f?-��q͏�D�f�9�nƱ����cw�Y���n��߀                                                                                    �����N�2p6��)��9Ny8��$�XC�    ���s]n���m����w�[}�����������]w�V��{���߀                                                                                    ��� R �QAJ�$��Q*) QAED��$�d �Q    ���wA`�,j�����[~���5°����]w�[��{���߀                                                                                    ������QO"�$��+��=OE|��*�D �Q    ���w_o���j�����[n����������]w�]��{���߀                                                                                    ���R �QQ�$���*JEQE@��*�D �Q    ���w]n���wn���w�[}�5����������g�ֻ�{���߀                                                                                    ���R ��QJ�$��P�)DEQED"�)D �S    ���wcq�.?�q�p͏�[~wv9�;°������ٺ�|r��߀                                                                                    �����H��2p������=Oy8h&E ��    ��������������������������������������߀                                                                                                    �                    ���������������������������������������߀                                                                                                                        ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ��������������������������������������߀                                                                                            �          @          ��������������������������������������߀                                                                                            �         @          ��������������������������������������߀                                                                                            �         @          ���8��ӎ9���c�Ɏ2'g���64����?����p��߀                                                                                   �,,q�8��p6q���+J��Nv8�s8<�    ����M�Muֻ��}mw�w����}���}�����������߀                                                                                    ���)D���$�)%P,�K*,�AIE 
DEQ    ����]��uۃ��am����}U��}�������.��߀                                                                                   �"�$|���$��%�P(��*�OI|�z|E�    ����]��uݿ��]m�}�����}U��}����u������߀                                                                                   �"�"@���$�)%P(��*�QI@@�@E    ����]�]uֻ��]mw�u����~���}����u�����߀                                                                                   (���)D���$�)%P(�*(�QIE �DEQ    ���8]�ݎ9���am�����~��7}���?����p��߀                                                                                   Ǣ"q�8��pq�$�H(�)ȂOI8�z8<�    ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ��������������������������������������߀                                                                                                  @     �         ���������������������������������������߀                                                                                                      @          ���������������������������������������߀                                                                                                      @          �����8�ƛs�Ӈ�i������̔8�N2�S��������߀                                                                                   8�9d�,x3�<�`08V3k���`�	+',      ������}�j��Mwۦ��o�_���}�ֿM��WM����߀                                                                                   D(�� ��$YE��YJJ(�J)@�	,��      ������}����]w�.���_��ݵ�}�ֿ]�WW�����߀                                                                                   D/�=��'�E�@�<Q"J/�J)@�
��"      �����������]w�����_������ֿ]�WW�����߀                                                                                   D(E��$E �DQJ(J)@�
��"      ������}��m�]wۮ��o�_���}�ֿ]��W]����߀                                                                                   D(�E���$QE��DQJJ(�J)@�H��      ����������]��n������δ8��:�]��X�����߀                                                                                   8
'=L�x#�<�b <Q1K�I�@�H�"      ���������������������������������������߀                                                                                                                       ���������������������������������������߀                                                                                                                        ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ��������������������_�����������������߀                                                                                                 �  �               �������������������������������������߀                                                                                                  �  �                �������������������������������������߀                                                                                                  �  �                ���8��p�q�?1��4L6?T��c�
s�?�10���L�m�߀                                                                                   �+3��l��8��˳����d��
�q��';�9�   ����S[�����n���յ��S]�]j���u��W[]5���߀                                                                                    ��QAI �EA*J* ����R �)(����   ����WX.���`�X?u��WA�A����}��P[Au���߀                                                                                   '���OH��A����J+ਾ�EH
 �)(����=   ����W[�����o��[�����W_�_����}��W�_u���߀                                                                                   (��QH@�A� JJ* ���%D
 �)(�$��E   ����W[�����n�뻾յ��W]�]j���u��W[]u���߀                                                                                   (��QQI �EDA*J* ����R
 �)(����E   ���8Wlp�p�?q��5�6?Wc�c���ߎ6���cv���߀                                                                                   Ǩ���D��8�C��K�����d�L
 q�/'$��=   ���������������������������������������߀                                                                                                                    ��������������������������������������߀                                                                                                      �          0   ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          �������o�������������������������������߀                                                                                        �       @ (                  �������_�������������������������������߀                                                                                        �      @ H    @     $   @     �������_�������������������������������߀                                                                                        �      @ H    @     $   @     ���8���O��q�8���18�N2��7}8ݏ�q�a�4��߀                                                                                   �'3 �$�@�8�X�i����`IȂ�"p5��i�    ����W[_��鮺�}����}�ֿ��|�]wٮ�����߀                                                                                   (����%AQE(�eH)(�J)@J(� ��&QQJ,�   ����W]�_�����p}���}�ֿ��}�k۠�����߀                                                                                   �� �%AQD��E�I�/�J)@J(�'��$_QJ(�   ����W^�_��������������ֿ��}�kۯ�����߀                                                                                   �� �%AQDHE J)(J)@J(�(��$PQJ(�   ����W[_��>뮺�}����}�ֿ��}�wwۮ�����߀                                                                                   (�����QE(�EJ)(�J)@2)�(��$QQJ(�   ���8���_����8������:��9}�w���a�7�߀                                                                                   �'# ��@�N8�D�I�'I�@!Ƃ'�pN�)Ȁ   ���������������������������������������߀                                                                                                                        �������������������������?�������������߀                                                                                         `                �              ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ��������������������������������������߀                                                                                     B  (            �                  ��������������������������������������߀                                                                                       H            �                 ��������������������������������������߀                                                                                       H            �                 ���3�8ϖ18�8����~8��c�3�㍌���������߀                                                                                   �Z�0i���'3 9��;<��r��Hrs0          ������_���}�W[���[]]mt���uu���������߀                                                                                   (S(�H)(�(���E(�����(H"��H          ������_��}�W]����[]Am���uu���������߀                                                                                   (R/�I�/��� E�����(�H ��           ������ߵ����W^����[]_m}���uu���������߀                                                                                   (R( J)(�� E�����)H ��          ������_���}�W[���[]]mu����uu���������߀                                                                                   (R(�J)(�(���E(�����)0"��H          ���7��߶��8�����8�Ccm���㍍���������߀                                                                                   �J' I�'�'#9�$���r$� rr2          ���������������������������������������߀                                                                                                                          ��������������������������?������������߀                                                                                                           �              ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          ���������������������������������������߀                                                                                                                          �                                      ����������������������������������������                                                                                   �����������������������������������������                                                                                                                           �����������������������������������������                                                                                                                           �����������������������������������������                                                                                                                           �����������������������������������������                                                                                                                           �����������������������������������������                                                                                                                           �����������������������������������������                                                                                                                           