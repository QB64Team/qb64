�i  ,|��                       �       0  0                                             �       0  0                                             �       0  0                                             �       0  0                                            3 � `                                                    3 � `                                                    3 � `                                                    3 � `                                                    0 � `                                                    0 � `                                                    0 � `                                                    0 � `                                                    0<�p<x�<7�                                           0<�p<x�<7�                                           0<�p<x�<7�                                           0<�p<x�<7�                                           fٳ`�6f�ـ                                          fٳ`�6f�ـ                                          fٳ`�6f�ـ                                          fٳ`�6f�ـ                                          ~߰`>��6~1��                                          ~߰`>��6~1��                                          ~߰`>��6~1��                                          ~߰`>��6~1��                                                                                                                                                              `�0`f��6`3                                                                                                                                                                                                                         3fٳ`f͛6f��                                                                                                                                                                                                                        <�0>x��<7�6�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��            ��            ��            ��                                                                                                                                                                                       �"|           �"|           �"|           �"|          ݀            ݀            ݀            ݀          "             "             "             "                                                                    �ǀ          �ǀ          �ǀ          �ǀ         � 8            � 8            � 8            � 8          D            D            D            D                                                                   8�$x�          8�$x�          8�$x�          8�$x�        ۇ           ۇ           ۇ           ۇ         $ �          $ �          $ �          $ �                                                                  ϟ�Ϙ          ϟ�Ϙ          ϟ�Ϙ          ϟ�Ϙ        0` 0`          0` 0`          0` 0`          0` 0`         � H            � H            � H            � H                                                                  |����         |����         |����         |����        �            �            �            �          D            D            D            D                                                                   ��$��        ��$��        ��$��        ��$��      8� �         8� �         8� �         8� �        $           $           $           $                                                                  ?O���@        ?O���@        ?O���@        ?O���@      �� h�        �� h�        �� h�        �� h�        H �            H �            H �            H �                                                                  o������        o������        o������        o������        @          @          @          @      !           !           !           !                                                                   �����|�        �����|�        �����|�        �����|�      &   �         &   �         &   �         &   �           @             @             @             @                                                                ?������       ?������       ?������       ?������      �`   0        �`   0        �`   0        �`   0           �             �             �             �                                                               �������       �������       �������       �������     1    d       1    d       1    d       1    d      ��           ��           ��           ��                                                                  �������       �������       �������       �������                                                @             @             @             @                                                                    �� ����      �������      �������      �������     � �          �             �             �                                                                                                              ��� �{@      ������{@      ������{@      ������{@    	 x � ��      	     ��      	     ��      	     ��         B            B            B            B                                                               -��  �ݠ      -������ݠ      -������ݠ      -������ݠ     �  "@            "@            "@            "@                                                                                                                        [��   ���      [��� ����      [��������      [��������    $@          $@ �         $@            $@                 @             @             @             @                                                              ��   ?��      ��� ���      ��������      ��������     �   �        � 8 �         �             �          @     �      @     �      @     �      @     �                                                              ���   ��      ���  ���      ��������      ���������    Q      P      Q �  P      Q  �  P      Q      P    �             �             �             �                                                                    o�    ��     o��   ���     o��� ���     o��������    � �    H      �     H      �  <�  H      �       H                                                                                                               ��    ��     ���   ��     ���  ���     ���������                �       �                                                                                                                                    ��    ��     ���   ?��     ���  ���     ��������   @          @    @      @          @  �                                                                                                              ��     �o     ���   �o     ���   ��o     ���� ?��o   H     �     H `   0 �     H     �     H  �  �    �             �             �             �                                                                    o�     �     o�    ��     o��   ?��     o��� ���   �     �@     � �    @     �    � @     �  ` 0  @                                                                                                                   
��     ?��    
��    ���    
���   ���    
���  ����        @                                  �               @             @             @             @                                                             ��     ?��    ��    ���    ���   ���    ���  ����        @                  @                                                                                                                                  ��     ��    ��    ���    ��    ���    ���   ���  
             
           
  �         
    �                                                                                                                    ��     ��    ��     ���    ��    ���    ���   ?���  
 @          
           
           
     @     @              @              @              @                                                                     =��     ��    =��     ��    =��    ���    =���   ���  @@      @    @     � @    @      @    @        @                                                                                                                  /      ��    /�     ?��    /�    ���    /��   ���  ��          �     @     �          �                                                                                                                          +�      ��    +��     ?��    +��     ���    +���   ���   �                @                  @        �              �              �              �                                                                     k~      ��    k�     ��    k�     ���    k�    ���  �            �             �           � �                                                                                                                            ^�      �p    ^��     �p    ^��     �p    ^��    ��p  !       �    !         �    !      � �    !  �     �                                                                                                                  W�      ��    W��     ��    W��     ��    W��    ���  (           (             (      �     (                                                                                                                         V�      ��    V��     ��    V��     ?��    V��    ���  )            ) @           )      @      )                                                                                                                              ~�      �P    ~��     �P    ~��     ?�P    ~��    ��P         �     @      �          @ �           �  (              (              (              (                                                                      ��      ��    ���     ��    ���     ?��    ���    ���  P           P @          P      @     P                                                                                                                         ��       ��    ��      ��    ���     ?��    ���    ���  R            R �           R      @      R                                                                                                                              ��       ��    ��      ��    ���     ��    ���     ���              �                                @              @              @              @                                                                      ��       ��    ��      ��    ���     ��    ���     ���  @      @    @ �     @    @        @    @      @                                                                                                                  ��       ��    ��      ��    ���     ��    ���     ���  R            R �           R              R                                                                                                                              ��       ��    ��      ��    ���     ��    ���     ���  R            R �           R              R                                                                                                                              ��       ��    ��      ��    ���     ��    ���     ���         P      �     P             P           P  R              R              R              R                                                                      ��       ��    ��      ��    ���     ��    ���     ���  R            R �           R              R                                                                                                                              ��       ��    ��      ��    ���     ��    ���     ���  R            R �           R              R                                                                                                                              ��       ��    ��      ��    ���     ��    ���     ���  @      @    @ �     @    @        @    @      @                                                                                                                  ��       ��    ��      ��    ���     ��    ���     ���              �                                @              @              @              @                                                                      ��       ��    ��      ��    ���     ?��    ���    ���  R            R �           R      @      R                                                                                                                              ��      ��    ���     ��    ���     ?��    ���    ���  P           P @          P      @     P                                                                                                                         ~�      �P    ~��     �P    ~��     ?�P    ~��    ��P         �     @      �          @ �           �  (              (              (              (                                                                      V�      ��    V��     ��    V��     ?��    V��    ���  )            ) @           )      @      )                                                                                                                              W�      ��    W��     ��    W��     ��    W��    ���  (           (             (      �     (                                                                                                                         ^�      �p    ^��     �p    ^��     �p    ^��    ��p  !       �    !         �    !      � �    !  �     �                                                                                                                  k~      ��    k�     ��    k�     ���    k�    ���  �            �             �           � �                                                                                                                            +�      ��    +��     ?��    +��     ���    +���   ���   �                @                  @        �              �              �              �                                                                     /      ��    /�     ?��    /�    ���    /��   ���  ��          �     @     �          �                                                                                                                          =��     ��    =��     ��    =��    ���    =���   ���  @@      @    @     � @    @      @    @        @                                                                                                                  ��     ��    ��     ���    ��    ���    ���   ?���  
 @          
           
           
     @     @              @              @              @                                                                     ��     ��    ��    ���    ��    ���    ���   ���  
             
           
  �         
    �                                                                                                                    ��     ?��    ��    ���    ���   ���    ���  ����        @                  @                                                                                                                                  
��     ?��    
��    ���    
���   ���    
���  ����       @@          @            @      �   @                                                                                                                       �     �     �    ��     ��   ?��     ��� ���   �     �      � �          �    �       �  ` 0                                                                                                                          ��     ��     ���   ��     ���   ���     ���� ?���                `   0                    �                                                                                                                         ��    ��     ���   ?��     ���  ���     ��������                  @                  �                                                                                                                         ��    ��     ���   ��     ���  ���     ���������                      �           �                                                                                                                                          ��    ��     ���   ���     ���� ���     ���������     �                       <�                                                                                                                                       ��   ��      ��  ���      �������      ��������    �             � �         �  �         �                                                                                                                               ���   ?�x      ���� ��x      ��������x      ��������x    @   ��      @ 8 � �      @     �      @     �                                                                                                                        o��   ���      o��� ����      o��������      o��������         @        �   @             @             @                                                                                                                        ?��  ���      ?��������      ?��������      ?��������      �                                                                                                                                                                         ��� ���      ��������      ��������      ��������     x � B            B            B            B                                                                                                                         ��� ����      ��������      ��������      ��������     �                                                                                                                                                           �������       �������       �������       �������      @             @             @             @                                                                                                                              �����       �����       �����       �����      ��           ��           ��           ��                                                                                                                            ������|       ������|       ������|       ������|           �             �             �             �                                                                                                                          �������        �������        �������        �������          @             @             @             @                                                                                                                           ]������        ]������        ]������        ]������      "           "           "           "                                                                                                                             ߷�o��        ߷�o��        ߷�o��        ߷�o��        H �            H �            H �            H �                                                                                                                            ������        ������        ������        ������       $           $           $           $                                                                                                                            �����         �����         �����         �����        D            D            D            D                                                                                                                              �o���          �o���          �o���          �o���         � H            � H            � H            � H                                                                                                                             7���`          7���`          7���`          7���`        $ �          $ �          $ �          $ �                                                                                                                            ����          ����          ����          ����         D            D            D            D                                                                                                                             ���           ���           ���           ���          "             "             "             "                                                                                                                               ��            ��            ��            ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           ?                        ?                                                                                                                                                                                                    0             3                          3                                                                                                                                                                                         0             0                          3                                                                                                                                                                                         >���          0���          ���          3���                                                                                                                                                                                      3훰          >훰          훰          훰                                                                                                                                                                                      ̓0          3̓0          ̓0          3̓0                                                                                                                                                                                      ̓0          3̓0          ̓0          3̓0                                                                                                                                                                                      3͛0          3͛0          ͛0          3͛0                                                                                                                                                                                      ��0          ��0          ��0          ��0                                                              