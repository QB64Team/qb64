�Vb  dN`r              x         l   �                           x         l   �                           x         l   �                           x         l   �                           � ��     �   �                           � ��     �   �                           � ��     �   �                           � ��     �   �                           � ��     �   �                           � ��     �   �                           � ��     �   �                           � ��     �   �                           ��<y����<���<�8                          ��<y����<���<�8                          ��<y����<���<�8                          ��<y����<���<�8                          y�f́���6f���3fٰ                          y�f́���6f���3fٰ                          y�f́���6f���3fٰ                          y�f́���6f���3fٰ                          �~�����6f�͘0fٰ                          �~�����6f�͘0fٰ                          �~�����6f�͘0fٰ                          �~�����6f�͘0fٰ                                                                                                                  �`�����6f�͘0fٰ                                                                                                                                                              ͛f́���6f�͘3fٰ                                                                                                                                                              x�<x�ٞ��<�͘<�3l                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            8                 �                8        |                �                |                                                                                                |                �                |        |                �                |                         @                                         @                       }                �               }       }                �               }       �                �               �       9                �               9       }                �               }       �                �               �       �               B               �                        @                       8�               �               8�      }�               �               }�       @                               @                                                  d L              �0               @      f �              �0               �                         �                                                                 � #                �              h ,     � c              0�              l l     �               � |                    �                                         �                            �       !�               �             � #     � �             �              �        �                            �       !�             |  ��              �     !�             |  ��              �    � �             � �            � �      �             |  �              �    g !�            �  �0             !�    g !�            �  �0             !�    � �            �� �            � �    g  �            �  0              �   � a�            0�            g !�   � a�            0�            g !�   �� �            �� �            � �   �  �                          g  �   � a��           0�           � a�   � a��           0�           � a�   � ��           �� �           �� �     ��                        �  �   � ���           ~8��          � a��  � ���           ~8��          � a��  � �0           a�� ��          � ��    �0           `   �            ��  � ���          �8��          � ���  � ���          �8��          � ���  `� �          ��� �0          � �0  `  �          �   0            �0 �� !��          �  ��          � ��� �� !��          �  ��          � ��� �� �          �� �          `� � �  �                        `  � ��  ���         �  �         �� !�� ��  ���         �  �         �� !��  � ��         �� ?�         �� �    � �                      �  � ��  ��0         7�8  ���        ��  �����  ��0         7�8  ���        ��  ��� � ��         8�  ��         � ��   � 0         0 8  ��           � �p��  ��         ��8� ��`        ��( )��0p��8 8��         ��8  ��`        ��( )��0? ~8 8��         ��� '��         � ��0    �          � 8  � `           � 0���� �        ��3� y��8        p��� ������ �        ��0  ��8        p��� �� x� <�        ��@ I��        ? ~` ��p               � 0  � 0        0    � p��P ��        �����8        ���T T��p��� ��        ��    �8        ���t \�� c� w��        ��� rx�         y� #<�p              �       8        p       p��H %#�        ��?� ���8        p��H %#�p��� ?��        ��    �8        p��� '#� x =��        �'  ���         f0 ��p  �           �       8        p       0�%( )H�        �������8        p��* �K�0�?� ���        ��    �8        p��: ���? =� �x�        � �� � �         � F0�0  �         �       8        p       0��� JR>        �������0        0��� JR�0��� �>        ��    �0        0��� Nr�? �� {��        �s�9��        ? c 1��0 @           �       0        0       �R� R��        ������|0        0�ҕR��������        ��     |0        0��s��������        �	�p�r�        ?�b �c� ! !         �       0        0�    �JR ��"         �?�����         �JR ������ ���         �               ��r ��{� ����         �'9�s���        1� c�� �  B          �                     � 5)K�)X          �������         ��K�/Z /�����          �@     D         ����?�=�{��x�         ���<��#�        �0 �1� � B�          �                �    ��))JZ          �����          ��( )K^  ������           �                ��99�~ ����{�          rs���9��        c� �1�� (B �(                            a      Z�� JR�          �����|         Z�� J^� ��� ���                 �         {�� �� ��� {��          A�s�9�p@        �c 1�b  )B �!(                            `      ZR� ��          ������          zҐ ��  o�� ��           @     @          ~� s��  {�� ��          9�p�s�          1�` c  ! aP                            0�     -JH $�h          ������          �zJ ��j  ��� ���                          ��z ��z  �{� ��           �9� ��          F1� C�  �0 BP                            0   @  -)$ I)h           �����`          =i$ I-x  7�� ��                 �          ?y� O=�  =�< y�x           ��<�           � 0�0  
� �                            @   0  �� RJ�          ������          V��Rz�  }����|                          ^��s��  w���{�           s�p�9�          #b �1�  
C !��                               0�  �R ���           o�����          �R ���  �� ���                          �r ���  �� ���           Ny�s�@          a� c`    a@                                `  IJ �%�           ������          +OJ���  >������                          /΂���  ;�{���           9�8��          �1�  0� B@                               �   5))Y�           7�����          5))Y�  ����`           @   B           �99��  =��y�           '���<�          � �0�  � ��                               �  ��JZ`           ?��߀          ��EK�@  ������            �               ��E���  ���{�`           >s�9π           c�1�   (B �)�                             c  �    Z��R�            ���|           Z��R�   �����                 �           {��s�   �����            �r	�p            �c�b    ) !(                                      ZR���            �����            {Ң��    o����             @   @            ��    {����            9�s�            1�Dc    !P                              1�     -JD�h            ����            �JD�j    �����                            ��D�z    �{ǽ�             �9��            F1��    � BP                                 @    -))h             ���`            =�/x    7����                 �            ?��?�    =��x             ���             � �0    
��                              � 0    �|J�            �����            V�|J�    }���|             �             ^����    w�|{�             s��9�            #|1�    
C���              �               | �    ���             o���            ��    ����                          ����    ���             N��@            a�`    ��@                            a�`    F(Š             �����            +F(Ũ    >�8��             �             /~8��    ;��Ǹ             9��            ���    > �@                             �     1�             7�@��            1�    �8?`             `��             �8?�    ���             '�_��            ���    �>�              `@�             0�    `l@             ��?�            `lP    �|�             ��0             �|�    ��p             ��             ��     � �             � 0              `      ��              �             ��     ��             �             ��    ��              ���             ��     ���             �             ��     ���             �             ���    ���             �             ���    ��߀             ��~             ��߀    ���                          ���      x               0�               x       x               0�               x     ���             ���             ���      `               0�               `     �               ` p             �      �               ` p             �      ���             ���             ���    �               ` @             �      p               �              p      p               �              p      ����             ���             ����    p                �               p       `�              !��             `�     `�              !�             `�     �}��             >���             �}��                      �                       ��              ?             ��     �D`             	�            �D`    ���             !���             ���    @                !                @       � �@            �             � �@    � P            �  @            � P    ����             s����            ����    �  @             r               �  @    �8B�            ��
�            �8B�    ��D�            ��            ��D�    k���            ����@            k���    b�               �                b�      �	�              �'��            �	�     � �            �           � �    ����            ����@            ����    �                                 �       ��0�            g           ��0�   �8�             @�C�           �8�    ����            ���@            ����    �                                 �       �0             d�@           �0    �Ơ            +�@            �Ơ   �u9_�            ����           �u9_�                                            ���            �HBC            ���    �� �            ��            �� �   �~T�             ��S�            �~T�                                             �|8o             E��            �|8o    ���            G��            ���    �|              �A�              �|                       D                       ��             �A�            ��    ���            ���            ���    ?T              �AP@             ?T                                                 ��D             ��             ��D    ����             ���            ����     }              p�@             }                                                 k��             ��Cx             k��     ��(�             ����             ��(�     �                \              �                                                  >w�              ��x             >w�     ��             ���             ��       �                �                �                                                   ��              ��              ��     >{��              ���             >{��      |@               �               |@                                                  ?��               ���              ?��      }�|              ���              }�|       �                               �                                                  }�               }��              }�      >��               ���              >��                                                                                        ��               >O�              ��      ��               ��              ��                        @                                                                   ��               �               ��      ��               ?��              ��                                                                                              �                �               �       ��               �               ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��  ��           � �           �    ?`                                                                                                                                     �  ` ��           � �           l    0                                                                                                                                      �  ` ��           � �               0                                                                                                                                      �y�s���|p         ��́�|p         ����0o�                                                                                                                                    ��fl��v�         �6o�v�         ٛm�>n�                                                                                                                                    �}�g���f`         ���f`         ٛm�0l�                                                                                                                                    �ͳf��f0         �6�f0         ٛm�0l�                                                                                                                                    �ͳfl��f�         �6m��f�         lٛm�0l�                                                                                                                                    �}�3���fp         �����fp         ���l�0l�                                                                                                                                                                                                                            