��`  Ta�                                                                         ������������������������������������                                                                                                            ������������������������������������                                    ������������������������������������                                    ������������������������������������                                    ������������������������������������                                    ������������������������������������                                     ?������������                 ���� ��           �����������������   � ?������������                 ����                                     ������������������������������������                                    ������������������������������������                                     ?������������                 ���� ��           �����������������   � ?������������                 ����                                     ������������������������������������  `  �                        pp  ������������������������������������  `  �                             ?������������                 ���� ��`      ����������������� 8�� ?������������                 ���   `                             ������������������������������������  <`                         �  ���������������������������������?��  <`                              ?������������                 ���� ��<|y���ϟp����������������� �� ?������������                 ���   <|y���ϟp                       ������������������������������������  ff͛�lٳ`                      ������������������������������������  ff͛�lٳ`                        ?������������                 ���� ��ff͛6lٿ`����������������� �� ?������������                 ���   ff͛6lٿ`                       ����2d��ɓ&O������������������������                                �  ���������������������������������?��                                     ?<�2D��ɓ&L��                 ���� ��           ����������������� 8�� ?������������                 ���                                     ��<��~�0`������������������������                                pp  ������������������������������������                                     ?������������                 ���� ��           �����������������   � ?������������                 ����                                     ������������������������������������                                    ������������������������������������                                     ?������������                 ���� ��           �����������������   � ?������������                 ����                                     ������������������������������������                                    ������������������������������������                                    ������������������������������������                                    ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            �����������������o�����������������                                                                                                            ����������������?�������������������                                                                                                            ����������������?�������������������                                                                                                            �����������1��?�Ɏ6��w������������                                                                                                            ����������2dɓ��?��u��[�������������                                                                                                            ����������2d���?��XX7������������                                                                                                            ����������2d����?��}�W[�������������                                                                                                            ����������2dɓ��?��u۷[�������������                                                                                                            �����������3���ێ;�\w������������                                                                                                            �����������|������������������������                                                                                                            �����������|�����������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                           ������������������������������������                                                              �                                             �����������}������������q�������                                                             @@                                             ��������������������������뮿������                                                             �                                              ��������������������������뮿������                                                             �                                              �����	�O�ߘ�M�|;_��a������뮇������                                                             �                                              ��������ؿ]5u�����n��o��ۮ�������                                                             �                                              �����녷�޸]u~��������������������                                                             �                                              ������u��޷]u}����������{��������                                                             @@                                             ������u��ܷ]uu���������������������                                                              �                                             ���������Cu�|=��a�q�*���q�������                                                                                                           ������������������������������������                                                                                                            �����������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ����������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ��������ޘ�1���8���18���ls�J�������                                                                                                            ����������]~��������v��髭�Z�������                                                                                                            ��������߷]p�������n�����Z�������                                                                                                            ��������߷]n���������������Z�������                                                                                                            ��������߷]n��������^�뫭�Z�?�����                                                                                                            ��������߸�p���8������s�j������                                                                                                            �����������������������������������                                                                                                            ��������������=���������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������?����������������                                                                                                            �����������������������������������                                                                                                            ������������������������������������                                                                                                            ����������ߍ8]���������������������                                                                                                            �������������]����?Z���������������                                                                                                            ����������߅�]�����n���������������                                                                                                            �����������u�]u�����v���������������                                                                                                            �����������u�Yu����Z���������������                                                                                                            �������������e���8f���������������                                                                                                            �����������������������������������                                                                                                            ���������������?��������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ��������������������������������                                                                                                            �����������������������u{�����������                                                                                                            �����������������������}�����������                                                                                                            �������������&�_���6��}�����������                                                                                                            �����������ߺ�������û������������                                                                                                            �����������ߺ�������ݻ������������                                                                                                            �����������ߺ�������݃������������                                                                                                            �����������޺�������}u{�����������                                                                                                            �����������������V7C}�������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            �����������������0�������������                                                                                                            �������������������]}��������������                                                                                                            �������������������_}��������������                                                                                                            ���������������_���_}����a�X������                                                                                                            ��������������m�����mm����]������                                                                                                            ��������������m����}}�m������߇����                                                                                                            ��������������mu���}}�ݭ�����w����                                                                                                            ��������������mu���]}��nm���]�w����                                                                                                            ��������������m�_�0�,����X�c�����                                                                                                            �����������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                    