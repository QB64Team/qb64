�[   ��F                                                                ������������������                              ������������������                                                                               ������������������                                               @                                               @                              ������������������                              ������������������                                                                                                                                ������������������                              ?������������������                              @                                               @                                               ?������������������                              |                p                              �������������������                              �������������������                              |                p                              �                 8                             ������������������                             ������������������                              �                 8                     8       �                           �                 ������������������                     8       ������������������          �                 �                                      |       �                           �                 ������������������                     |       ������������������          �                 �                                      �       �                           �      �        #�������������������        �         �       #�������������������         �      �        �                          �         �       �                 �         �      � (�      C������������������@       D         �       C������������������@         p      � 8�      �                 �       �     �  �       |                 �      |  �      ��       �������������������          �     �  �        �������������������       |  �      ��      |                 �         �     �  �       >�����w�������?�����      �  �      ��      A �� �    ?� �       0      �  �       A���p ����� ?��      �  �      ��      >�����w�������?�����       0      ?�  ~       }�����������߇��~{�p     �  �      ��      � � � �    �~��       0      ?�  ~       ���������߇� x?�     �  �      ��      }�����������߇��~{�p       0      � 8       ��?���� |9���q�=���8     ��@�      �C�      �         p����       8b     � 8      ?� �� |9����< <�     ��@�      �C�      ��?���� |9���q�=���8       8b     �        �������������������     ���       ���       �  ��    � ����       8D     ~�         � ��� ���� �� �     ���       ���     �������������������      (8D     �  �    ��������������      ��@      ��	�     @ �  ��   � ���     @<H     x�  �    _�� �� ���� � �     ǀ@      ��	�     ��������������      x<H     ��x���    �y�������}��������     ��ǯ ?�    �
�      �x�  ��   � ����      <8P�    ��x���     �����  }��� � ���    ǃǯ ?�   ���     �y�������}��������      8?���    �y���    ��~������������?=����    ��Ϯ �    �
?�     A ~�  ���  � ���@      <0Q��    �y���    A� ����  ��� ?< ��@    ��Ϯ �    ����     ��~������������?=����      ����    ?�`
��    }�~������������������    �C V ��   @�?�     � ~�  ��� ������� �      �0i�    ?�`��     �� ����  �  > ��     �C  ��   @���    }�~��������� �������     �0?�    �  �    >���?��������=�8���     �� � ��   ��?�@    A     ��� ��8  �     ~0��    �   |    A��?��  p   < �     ��   ��   �?�?��    >���?�����p  =�8���    �0	�    �  �    }���������������{����@p     |  @ ��  ��	�     ��     ����  ~�   �    �~pH�	    �   <    �������      x���?�     |    ��  ����    }�����������    {����@p    �~p�     p  �    ����0����������������`8      �  ��  	����  � 0   ���   ��   �    O�|p��     p  <   � ����       |����      �  ��  	�����   ����0�������    }����`8    O�|p��    � ��   �����}�����������o� ?�      � ��  ����    ?��   ��� � ``   �    o�8<�    �  �    � }���       � ?��      �  ��  ���"    �����}������    o� ?�    o�8<�q     � ��   �����������������  �      � �  ��&r�    ���  ����� 1���    /�93���      �  �   @� =���       �1����      �  �  ��r    �����������    �1���    /�83���      � ��   �����������������   �      � ?� ��g*?�     ����  ����  | �����  ��81Q�       �  G�    � � ���       �������     � ?� ��g*<@    ����������     �����   ��81Q�       p ��   ���o��������������   |�     � � ��7�$o�    A����  ��    ����@  ���q#       p  ��   A  ` ���        ����}�@     � � ��7�&l�   ���o�������  @   ����|�  ���q3g �  8 � �   }��o��������������   ?�  �    �  �?�gO��    �����  ��    �������    ?���:~7   8     @    �  ` ���        }�����   �     �  �<~gNF�   }��o�������      }�����   ?���:r7�  | �   <   >���o��?����������    �  � >   �  ��G��   A����  ��0    `A����   ���<pn   |      <   A  ` ?��        =����  �     �  �>G��   >���o��?���  �   =���� �   ���<po�  | �      }������������������   �p  �     x  ��F�3�   ����� ���    !����?�   ���4a�   l        �  � ��         ������  `     x  �F�3�   }��������         �����p   ����4a�x  �8�  ǀ  ������������������   �8  ��   <  ������   ����        !�����   �����   � �  ǀ  � �          ������  �    <  ��ҟ����  ��������          �����8  >����<  �|�  � ���?���������������   �  ��     ���t��   #� �� x       �����   �����`   �    � 0 ?� ��         ������  �      ���t��� ���?�����         �����  ����` �|�  �  �����������������   �  �>   ?�  ����	O� A� ����     �����   ���#�J~ �    �  x��           ������   �    ?� ��?�	O� ������          �����  ���#�J~   |�  �� �~����������������   �   �   ?� ������ `  �  ����     ������ ����/�@        p�  ��� =�          ������        ;� ������� �~�����          ����  ���/�D �8    �� ����y�{������������   ~� �    ?�  �����L  A   �          B����@  ǿ�?��` �     �� A���x {�          ����@       ?� ������L� ����y�{�         ���~� ~��?��g      �p }C� x��������������  � 8    p � �����   �  �x `�         !?��� �   ������       �p  �C�� ��           �����  8      ������p }C��x��         ����� 8�������     �p >��� ���������������  ��� 8    � � �����?� A  ��  �          0����   ?�������       �p A�����            _���� 8      ������?� >������           _��￀� 8?�������      8 }��~ ��������������  ��p p   p�  � �������� �  ��          G��  ?� ������       8 ��~���           '����� p   p   �����d���� }��~���            '����p w����'.���     8 ����  ���������������  ���8 p   ��  !� ���`��   ��          @�   � ��� ���       8������           8� ���� p   �   !��{�` ��8 ��������        @   8� ���8 w��� ���  �?�  ����  ~�������������� ���� � �p  p� �_D�?�   ��         >       � ��� |�    �?�  ?����~�        >    ����� � �   p��D�?�������~�             ���� ���� � � �?� p���  }������������������� � �� � � ��J�  @ �� @       >      �  ��S���     ?�  ����}�        >   ������ �  �    ��J� �����}�       @    ����� �}�:S��x � �?� � ���  =������������������� � �� � � ��D���  � ���0�     >      �� ��#����  ?�    �������        >   �������� A�    ��D���������            ����� ��:#��?��<� � ����  =���������������  ~��@�� � � ��`��� A  ���!        >      �� ����� < @    A�������        >   �  ~����@ �   �<�G`�#��������� @          �  ~��;����  � � }���  ������������������   �p � p��p?�����  ���C        >  � ��� ���������    �  p ������݀        >    �  ��   p � p���p?�s��}�����݀             �����;�����p8 �  � y���  ��������������������� �  � p���r�a����  ���B        >   `���� x������� 8 H     ������݀        >    |  ���� @    p��Gr��#��y�����݀             }�������;���p8 �   � v���  �������������������� �  � 0�?��3������  ����        >   c��� 8����������8        �������         >      �8��        0�?�3����v������             �������y���?��8  �  p n���  ���������������������    � 0 =�_#����   ����           ��� ������ @8  �     �������               �؁�       08=�#���n������            �����	�����| px    �� _��  �����������������    t|  8@!�"p�	�   ���            ��� ������ H8     �� �����                  ���    |  0x!�"qp�_����     � �    ����������� xx   �� ?��?� ��������������������    .�  x@�� ��   ���            ��� �� ��� ��8   �� ���?���                  ���    �  px�� �?��?���       �    ��������� ��xx    �� ��� �����������������{��p   �  x@���@���    ��             ������ ��: �8    �� �����                  x��p   �  px���@������       	�    ���{����: �xx p  � ������������ ���������w�� � �� x@���� a�    ��            C����� ���� 8    � ������                  p��    �� px���� o�����       �    ���w����x�!x�  �  �� ��� ��~��������hW��������w�� � �� x�;����� !��      �             !����������D 8     �� ��� ��~                  p��    �� p�;���� /��� ��~       ��8    ���w����?��D x� �  �� ����������������������o�� � �� ��_���� ��� �              ��������� < <     �� ���  �                  `��    �� ��_�S��������       �|   ��o������8< �� � �� �x����������������������o�� ���� ������@`�� ��� @           ����� ������      �� ���  �                  `��   �� ���#��@`�x������      ��   ��o������ �� ��> �� ����������������������o������ �����  0�� ���             ���� 8��� � �   �� ��  �                  `��   �� ��S�� 0������        ��   ?��o��8��8�����>�� �����������������������o������� ��������� ���`x             ?���� p��XD?��  �� ���  �                  `��� @�� �������������       i�  � ��o��p>NHD?����p>� 9�߿��������������?�������o�����;����G�7O��� ?�����            /�����r?��|@��  � >�߀                      `�p� �����G�H�?�߿���         i�    ��o��r<x�D@���� ?� 9����������������?����������� �� ���� �� ?���              ��������X �@�  ?� >��                      ��p� @� ����	 ?�����         i�     �������XH �A�� �   � q�������������������������    � ���� �� ��� �           ������A �@ �   � ~��                     ��8    � ���� �����        9�    ������A �C��     � q���������������D}����������     | ����0�� ���8              ����w�A��      � ~��                    ���8     | ����0�����        ��    ������A��#���       ���������������D}���������       ����� �� ���@            @  � � ��� w��G�� �       ���                    ���       ������� ������         ���  ����� w��G�����       ���������������d��������7�       ����� �� ����               �   8�� G��G�  �       ���                    ���       ������� ������         �     ��7� G��G� ���     Ç��������������$�����������       ��r� �� ���              D   �� ��@�� �      ���                    ���Ȁ       ����r������          �    ����� ��@�����      ����������������$�����������       ��?
� �� ���                D   �� 9�P��  �      ���                    �����       ����?
������           �  @ @����� 9�P����  �   ����������������������������     <�� � ��               D   �� 8S��  �  �   ���                    ������     ?��������          ^     ������8S��?�� �   ��������������������� ��� �   x8� H� � ��                "   ��  0G�8 8 x �   ���                    � ��� �   �� J�����          Z     � ��� 0W�8�� �   <���������������������  7�� �  �8� M� � ��                "   ��   o� 8  �   ?���                    ���8� � �  ��� M�?����          z�    ���7��  o�	��� �   |��������������������   �� �  �8� BM�  � ���`                "   ��  "n  8  �   ���                     ��Ȁ � �  ��� BM� �����         c��     ����� "n��?���   � ��������������$�����   �� �  �p?�  �  � ���@                "   ���   ,  p ��   ���                    ����� | �  ��?�� � �� ���          ��@   ������   ,��?���  ���������������� o����   �� �  �p?�    � ����                !   ���   (  p ��  ����                     ����� > �  ��?�� ������           ߐ �   ������   (��?�� �  �����������������������   �π   > p?�  B  � ���                   ��� 0 "  p � �  ����                     ����� ?�   ?��?�� B������                �������0 "?���|     ���������������������    ���    � ��  �  � ��           ��      ���   $  � �    ����                     ����� �    �� �� �����           5    ���� ���  $����>    > <|��������������������    ���   ���     <� ?��            `       ���   8 � �    ?����                    ����� �   �� ��  ?��|��           �      ���� ���  8�����   � <���������������ʟ�����    ���   ���      <���               ���   0  � ��   �����                    ����� �   �� ���  ������          5`     ���� ���  0�����  � x���������������o�����    ��  � ��       x���          	       ��      �  ��  �����                    ����� ��  ��� ���  ������           T�     ���� ���  �������  ��x��������������j������    ��  ����    �x���          `�     ��     �  ?�  �?���                    ����� ��  ��� ���  ������  �        8�      ���� ���  �������� ���������������j������    ��� �x���     ��� �          	      ���    x�  ����� ��                    �����  ?� ��� �����������   �        �     ���� ��� ���������> ����������������������    ?����������    > ��� |          " ��      �?��   ��  A������ ��                    ����� ����� �����������x           U      ���� ?����������ǃ���������������������������    ?�<�����ǀ   ���� <           $@D�      �?�<   ��  8���� � ��                   ����� ������ ������������                  ���� ?������������  �����������������������    ��  �  ���  ����           D�"D      ���  �    ���?� � �                   �����  ����� �����������                  ���� �������� ���� �����������������������    ��� � > ���� ����@          I D      ���� � >   �?� �� � �                   �����  |���� ������������                 ���� �������� ����� �����������������������    ����  ~ ����� ����H         @I@  !   �����  ~   �  �� � �                   �����  ?�  ��� ������������                  ���� ��������  �� ?�  �����������������������    ����  �  �� ?�  ����@          ID   "   �����  �   ����� �  �                  �����  � ��   ������������                 ���� ��������  �     ? ���������������������    ��    �  �     ? ����         L�&H   "   ���    �   ������ �  `                  �����  �����   ������� ��`                 ���� ��������  ?��    � ���������������������    ��    �  ?��    � ����          $DD�   "   ���    �    ����  �  `                  �����  �����   ?������� ��`                  ���� ��������  ?��   � ���������������������    ��    �  ?��   � ����        " ��   "   ���    �    ?����  �  `                  �����  �����   ?������� ��`                  ���� ��������  ��   � ���������������������     ���   ?�  ��   � ����          	   D   � ���   ?�    ����  �  `                  �����   ����   ������� ��`                  ����  ��������  ��   � ���������������������     ��   �  ��   � ���1�          �3    D   � ��   �    ����  �  @                  �����   ?����   ������� ��@                  ����  �������  ��   � ����������������������     ?��  ��  ��   � ���!           `�    D   � ?��  ��     ����  �  �                  �����   ���    ������� ���                  ����  ?�������  ��� �� ����������������������     ��  �   ��� �� ���!               �   � ��  �      ��   �  �                  �����    ���    ������� ���                  ����  ������    ��� ?�� ����������������������     �����    ��� ?�� ���!            �`�   �   � �����      ��   � �                  �����    �      ������� ���                  ����  ������    �����  ����������������������     ������    �����  ���!            ?�      � ������            � �                  �����            �����  ���                  ����  ������    �����  ����������������������      ������    �����  ���!                    �  ������            � �                  ?����            �����  ���                  ?���   ������    �����  �~��������������������     �����    �����  �� a                   �  �����            � ~                   �����            �����  �~@                  ����   �����    �����  �����������������������     ����     �����  ���                <   �  ����             ��                   �����            �����  ���                  ����   ����      �����  ����������������������     ����      �����  � �                 >   �  ����             ��                    ����             �����  ��                  ���   ����      ���   p������������������������     ����      ���   � �                 ~   �   ����             ���                    ����             ���   p���                  >���    ����      ���   �������������������������    ��       ���   � �  @              �   �   ��              ���                   ����             ���   ���                  ���    ��        ?�    ��������������������������    ��        ?�    � �                 �   �   ��              ���                   c�����              ?�    ���                  c����    ��              �����������������������?�                     � ?�                !   �                    ���                   ��?��                    ���                  ��?�                     ��������������������������                     � ?��               B ���                    ���                   ����                    ���                  �����                       �������������������}��                    �������                �������               �����                   | ������                    �                 }��                    ������������������������{�m�����                   ��       �      �     �                             |       x b     �              ������        �       {�m�����               �������������������������7��������                  ���       �     ��     @                                    � 2     @              �������        �       ���������              ������������������������7��������                   ��@       ��     ��                                    �      �                     �������        ��      ���������              >    �����������?�������/���   �              A�������@       �@     `��?����              A�����          �      � ?����              >    ��        ��      ����   �              |    ������������������/���   �              ��������@       �      `���?����              ������          �      � ?����              |    ��        ��      ����   �              �    �����������|������ _���    �             �������        ~     � ��?����             �����          �      �@ ?����              �    ��        �      �_���    �             �    ����������������� _���    |             	�������        	�      ��?�����             	�����          |�     �@ ?�����             �    ��        ��     �_���    |             �    ����������ǔ������� _���    >             �������@       ��    8 ��?�����                 "          @      �@     �             �?�����        ��      �_�������>             �    ����������ϔ������ ����                 #�������@       �@   �0 ��?������            "    "           �     �     ��            �?�����        ��     ��������             �    �����������������������    �            G�������        �   � � ��?�����@            D    "          �     ��     �@            �m�۝��        ��     ������m���            p    �����������|�����������    �             ��������        ~    � ��?�����              �    "          �     ��      �             p?�����        �     �����������            >�    �����������������������    �            A�������      	�    ?� ��?�����            A    "          |�     �� 6     |            >�?�����        ��    �����������            }�    ���������������������a�    �            �?�������             �� �?�����            �     "                  � n     >            }�m�۝��    ����������?���m��m���            ��    �����������������������     �           �������             ?�� �?�����           @    "                  �� �                 ��?�����    ��������������������� �           �     �������         �������     |           ��������             ��  �?������           �    "      ���������  ���     �           � ?�����    ?��������������������� |           �     ������� 0 �  `������     >           ��������    0 �  `��   ?������                "      ��������  ���     �           ��I$]��    ?����������������$�Ih>           �     ������� 0?�`�������                #���������    0?�`��   ?�������          "     "      ��������  ����     ��          ���   ���    ?�����������������   ?�           �           8  A �  �     �     �          G�������������  ? ��  ������?������@          D     #���������������������     �@          ���   �      ?���������     �   ?��          p     ������8 � G�  ��������     �           �������     �   @8         ?������            �           ������7��             �           u��I$_������?�����������������$�Im�          >�     ������8 �  #�  ��������     �          A������     �              ?������          A           ��������             |          >���   �������?�����������������   ?���          }�     ������8   @    ��������     �          �?������     �   @           ?������          �            ����������             >          }���   �������?�����������������   ?���          ��            8 �@ �  �             �         ������������� �@ �  �������������         @     ?���������������������               ����I$@      ?����������      $�Im��         �             8 � 	  �             |         �������������� �� �  ��������������         �     ?����������������������     �         ���   �      ?��������         ?��|         �             8 �����  �             >         ��������������  ���  ��������������               ?���������������������     �         ����   �      ?����������         ?��>         �             8 �  	�  �                      #��������������  ���  ���������������        "      ?���������������������     ��        �m��I$@      ?����������      $�Im�         �             8   ���   �             �        G��������������   ���   ��������������@        D             ���  ���             �@        ����   ����   ?����������  ����   ?���        p             8 �����  �             �         ��������������� �����  ��������������          �             ��  ��              �         w���   ����   ?����������  ����   ?���        >�             8 � 	  �             �        A�������������� �� �  ��������������        A             ��������              |        >�m��I$m��nI$�?��������I$���m�$�Im���        }�             8 � 	�  �             �        �?��������������  �   ��������������        �              ������              >        }����   ����   ?����������  ����   ?����        ��             8 �@ �  �              �       ��������������  @   ��������������       @             �������                      �����   ����   ?����������  ����   ?����       �              8   @    �              |       ���������������   @    ���������������       �             ���������              �       �[m��I$m��nI$�?����������I$���m�$�Im��|       �              8 �  #�  �              >       ��������������� �  !�  ���������������                     �������              �       �����   ����   ?����������  ����   ?���>       �              8  D  �                     #���������������  � C�  ����������������      "              ���������              ��      �����   ����   ?��������  ����   ?���       �              8  � ��  �              �      G���������������   �0  ���������������@      D              �����x/��              �@      ��m��I$m��nI$�?����������I$���m�$�Im���      p              ; 0>�`�              �       ���������������� 0 ``���������������        �              ������_��               �       w����   ����   ?����������  ����   ?����      >�              ; 0 �  `�              �      A��������������� 0 �  `���������������      A              ��������               |      >�����   ����   ?����������  ����   ?����      }�              8         �              �      �?���������������         ���������������      �               ���������               >      }��m��I$m��nI$�?����������I$���m�$�Im�ہ�      ��              ?����������               �     ���������������         ���������������     @                                             ������   ����   ?����������  ����   ?��� �     �               ?����������               |     ����������������         ����������������     �                                       �     �����   ����   ?����������  ����   ?��� |     �               0         �               >     �����������������������������������������                    ���������               �     �F�m��I$m��nI$�0         �I$���m�$�Im�ې>     �                   $    `                    #�������������������������������������������    "               ����������              ��    �����   ����       $    `  ����   ?���      �                    �                   �    G������������������������������������������@    D        ?������������������������       �@    �����   �           �             ?��� �    p        ������    !�    ?�������        �     ����������      �����������      ?���������      �               ����������               �     rF�m��I$_������    !�    ?�������$�Im�ے�    >�        ������    �    ?�������        �    A���������      �����������      ?���������    A               ����������               |    >�����   �������    �    ?�������   ?��� �    }�        ������    O��   ?�������        �    �?���������      �����������      ?���������    �                ���������               >    }�����   �������    O��   ?�������   ?��� �    ��                  �@         �         �   �������������������������������?���������   @        #����������������������             ���$�Im�ۜ          ��         ��m��I$m��   �                   �@         �         |   ��������������������������������?����������   �        #����������������������         �   ��   ?���          ��         �����   ��|   �                   >|`         �         >   ���������������������~?����������?����������            #����������������������         �   ���   ?���          >�         �����   ��>   �                  �@        �            #�����������������   �    ������?�����������  "         #�������    |�   ������         ��  �m�$�Im�ۜ          ��         ��m��I$m�   �               B   ��       �         �  G����������������    ��   ������?����������@  D         #������    @   ������         �@  ���   ?���          ��         �����   ���  p               B   �@       �         �   �����������������    �@    ������?����������    �         #������     �    ������          �   w��   ?���          ��         �����   ���  >�               !   �@       �         �  A���������������    �     ���?����������  A         #�����    �    ���          |  >�m�$�Im�ۜ          ��         ��m��I$m���  }�               !   |@       �         �  �?����������� ��    ~     ?���?����������  �          #� ��    �    ?���          >  }���   ?���          �         �����   ����  ��               !   	�@       �          � ����������� ?��    	�     ���?���������� @         "� ?��    |�    ���            ����   ?���          ��         �����   ���� �          ��    ?����������     �          | ������������� � �  ��   ��?����������� �         "|7�����   @   ������          � �[m�$�Im�۝�����?�   ��   ���=���m��I$m��| �                ���������     �          > ������������������  �@  ������?�����������           #�������    �   ������          � ����   ?���     �   ��        �����   ���> �          �����p���������q����           #�����������8  �@  �   � � �?������������"          "8  ��   �   � � �          ������   ?��������w�   ��   q��������   ��� �          �����p����~����q����          �G�����������8  �@  {    � � �?�����������@D          "8  ��   �   � � �          �@��m�$�Im�۝�����w�   �   q�����m��I$m���p               p���������p    �          � ������������������   	�    ������?�����������  �          #�������   ~�   ������           � w���   ?���     w�   ��   p    �����   ����>�               p����������p    �          �A�����������������0  ��  @������?�����������A          #�������        ������           |>����   ?���     w�   ��   p    �����   �����}�               p���������p    �          ��?����������������� �   �������?������������           #�������   �   ?������           >}��m�$�Im�ۜ     s�   ��   ?p    ��m��I$m��A�{�               p���������p    �           �������������������  �    �������?������������@          #�������   �   ?������           {����   ?���     s�   ��   ?p    �����   �����w                p9����~���p    �           p�������������������  {   A ������?��������������          #������8   �   ������           �w���   ?���     p8   �   p    �����   ����pv                s����������p    �           p��������������������  ��  � ������?�������������           #�������   ~@   ������           �v��m�$�Im�ۜ     s�   ��   p    ��m��I$m��hpt                s����������p    �           p������������������� A  �@  ������?�������������           #�������   �  �������           �u����   ?���     s�  ��  �p    �����   ����pp                s����������p    �           p������������������� @� �   ������?�������������           #�������  �  �������           �s����   ?���     s�  ��  �p    �����   ����pp                s����������p    �           p�������������������  @ �   ������?�������������           #��������  �  Ϗ�����            �q��m�$�Im�ۜ     s��  ��  �p    ��m��I$m��npp                s�����~����p    �           p�������������     � 0 s  6 �    ?�������������           "     ���  �  �                �s����   ?���     s��  �  �p    �����   ����pp                r>���������|p    �           p�������������     �> ��  _ �    ?�������������           "     � �  ~@  |�                �s����   ?���     r>�  ��  |p    �����   ����pp                q��������p    �           p�������������     �� �@ �� �    ?�������������           "     � |   �  B�                �q��m�$�Im�ۜ     q�|  ��  ^p    ��m��I$m��npp                s����������p    �           p�������������     ��� �  �    ?�������������           "     � >  �  ���                �s����   ?���     s��  ��  ��p    �����   ����pp                s����������p    �           p�������������     ������   �    ?�������������           "     � ?  � ���                �s����   ?���     s��  �� ��p    �����   ����pp                s�����|����p    �           p�������������     ���0 �  �    ?�������������           "     � � � ���                �q��m�$�Im�ۜ     s��� � ��p    ��m��I$m��npp                s���������p    �           p�������������     ������   �    ?�������������           "     �  |@ � �                �s����   ?���     s�� �� �p    �����   ����pp                s��������|�p    �           p�������������     ���� �@ � ��    ?�������������           "     �   � 3| �                �s����   ?���     s��� �� 7|�p    �����   ����pp                s��������{�p    �           p�������������     ������ ��    ?�������������           "     �  � �x �                �vI$�F�m��I$\     s��� �� �{�p    �$�Im�ےI$�pp                s����������p    �           p�������������     ����� ���    ?�������������           "     � ���� �                �t   ����   �     s���������p    �   ?���   pp                s�����_����p    �           p�������������     �����  ��    ?�������������           "     � � ���� �                �t   ����   �     s���������p    �   ?���   pp                s���������p    �           p�������������     ���� ��  ��    ?�������������           "     � � ?�� �                �vI$�F�m��I$\     s���������p    �$�Im�ےI$�pp                s��|?���p    �           p�������������     ��� �� ?���    ?�������������           "     � �� � �                �t   ����   �     s�����?���p    �   ?���   pp                s���s����p    �           p�������������     ��� ������    ?�������������           "     � ��� � �                �t   ����   �     s����������p    �   ?���   pp                s���ߌ�����p    �           p�������������     ��� ������    ?�������������           "     � ?��� � �                �vI$�F�m��I$\     s���ߜ�����p    �$�Im�ےI$�pp                q���ߐ _����p    �           p�������������     ��� � _����    ?�������������           "     � ?��  @ � �                �t   ����   �     q���ߐ _����p    �   ?���   pp                r��ߠ _����p    �           p�������������     �� <� _����    ?�������������           "     � ���  � �                �t   ����   �     r��߸�����p    �   ?���   pp                s|���������p    �           p�������������     �| >?������    ?�������������           "     � ����   � �                �vI$�F�m��I$\     s|����������p    �$�Im�ےI$�pp                s��������w�p    �           p�������������     �  ������    ?�������������           "     �����     p �                �t   ����   �     s��������w�p    �   ?���   pp                s��������{�p    �           p�������������     �   ������    ?�������������           "     �����    x �                �t   ����   �     s��������{�p    �   ?���   pp                p��������p    �           p�������������     �  ��������    ?�������������           "     � �    8 �                �vI$�F�m��I$\     p��������p    �$�Im�ےI$�pp                s����������p    �           p�������������     �������������    ?�������������           "     �<      8 �                �t   ����   �     s�����������p    �   ?���   pp                s��������{�p    �           p�������������     ������������    ?�������������           "     �      x �                �t   ����   �     s���������{�p    �   ?���   pp                s���������p    �           p�������������     ����������{��    ?�������������           "     �          �                �vI$�F�m��I$\     s���������3�p    �$�Im�ےI$�pp                s��������p    �           p�������������     ���������y��    ?�������������           "     �           �                �t   ����   �     s��������y�p    �   ?���   pp                p��� ?�� �p    �           p�������������     �_����?�����    ?�������������           "     �           �                �t   ����   �     p_���� ?����p    �   ?���   pp                p��   �� ?p    �           p�������������     ����� �����?�    ?�������������           "     �           �                �vI$�F�m��I$\     q���� $����?p    �$�Im�ےI$�pp                p?��   ��  p    �           p�������������     �������������    ?�������������           "     �           �                �t   ����   �     s����  ����p    �   ?���   pp                p?��       p    �           p�������������     �����������    ?�������������           "     �           �                �t   ����   �     s����   ��p    �   ?���   pp                p��        p    �           p�������������     ������������    ?�������������           "     �           �                �vI$�F�m��I$\     r_��F��v�I$p    �$�Im�ےI$�pp                p��        p    �           p�������������     �������������    ?�������������           "     �           �                �t   ����   �     p������   p    �   ?���   pp                p��        p    �           p�������������     �������������    ?�������������           "     �           �                �t   ����   �     p������   p    �   ?���   pp                p �        p    �           p�������������     ������������    ?�������������           "     �           �                �vI$�F�m��I$\     rH�F��v�I$p    �$�Im�ےI$�pp                p           p    �           p�������������     ������������    ?�������������           "     �           �                �t   ����   �     p   ����   p    �   ?���   pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �t   ����   �     p   ����   p    �   ?���   pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �vI$�F�m��I$\     rI$�F��v�I$p    �$�Im�ےI$�pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �t   ����   �     p   ����   p    �   ?���   pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �t   ����   �     p   ����   p    �   ?���   pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �q��m�$�Im�ۜ     rI$�F��v�I$p    ��m��I$m��npp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �s����   ?���     p   ����   p    �����   ����pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �s����   ?���     p   ����   p    �����   ����pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �q��m�$�Im�ۜ     rI$�F��v�I$p    ��m��I$m��npp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �s����   ?���     p   ����   p    �����   ����pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �s����   ?���     p   ����   p    �����   ����pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �q��m�$�Im�ۜ     t�I$���m�$�Ip    ��m��I$m��npp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �s����   ?���     p   ����   p    �����   ����pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �s����   ?���     p   ����   p    �����   ����pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �q��m�$�Im�ۜ     t�I$���m�$�Ip    ��m��I$m��npp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �s����   ?���     p   ����  p    �����   ����pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �s����   ?���     p   ����  p    �����   ����pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �q��m�$�Im�ۜ     t�I$���m�$�Hp    ��m��I$m��npp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �s����   ?���     p   ����  p    �����   ����pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �s����   ?���     p   ����  p    �����   ����pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �q��m�$�Im�ۜ     t�I$���m�$�Hp    ��m��I$m��npp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �s����   ?���     p   ����  p    �����   ����pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �s����   ?���     p   ����  p    �����   ����pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �q��m�$�Im�ۜ     t�I$���m�$�Hp    ��m��I$m��npp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �s����   ?���     p   ����  p    �����   ����pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �s����   ?���     p   ����  p    �����   ����pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �q��m�$�Im�ۜ     sm��rI$�6�m�p    ��m��I$m��npp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �s����   ?���     w����   ���p    �����   ����pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �s����   ?���     w����   ���p    �����   ����pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �q��m�$�Im�ۜ     sm��rI$�6�m�p    ��m��I$m��npp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �s����   ?���     w����   ���p    �����   ����pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �s����   ?���     w����   ���p    �����   ����pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �q��m�$�Im�ۜ     sm��rI$�6�m�p    ��m��I$m��npp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �s����   ?���     w����   ���p    �����   ����pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �s����   ?���     w����   ���p    �����   ����pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �vI$�F�m��I$\     sm��rI$�6�m�p    �$�Im�ےI$�pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �t   ����   �     w����   ���p    �   ?���   pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �t   ����   �     w����   ���p    �   ?���   pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �vI$�F�m��I$\     sm��rI$�6�m�p    �$�Im�ےI$�pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �t   ����   �     w����   ���p    �   ?���   pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �t   ����   �     w����   ���p    �   ?���   pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �vI$�F�m��I$\     sm��rI$�6�m�p    �$�Im�ےI$�pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �t   ����   �     w����   ���p    �   ?���   pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �t   ����   �     w����   ���p    �   ?���   pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �vI$�F�m��I$\     sm��rI$�6�m�p    �$�Im�ےI$�pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �t   ����   �     w����   ���p    �   ?���   pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �t   ����   �     w����   ���p    �   ?���   pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �vI$�F�m��I$\     sm��rI$�6�m�p    �$�Im�ےI$�pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �t   ����   �     w����   ���p    �   ?���   pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �t   ����   �     w����   ���p    �   ?���   pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �vI$�F�m��I$\     sm��rI$�6�m�p    �$�Im�ےI$�pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �t   ����   �     w����   ���p    �   ?���   pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �t   ����   �     w����   ���p    �   ?���   pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �vI$�F�m��I$\     sm��rI$�6�m�p    �$�Im�ےI$�pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �t   ����   �     w����   ���p    �   ?���   pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �t   ����   �     w����   ���p    �   ?���   pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �vI$�F�m��I$\     t�I$���m�$�Hp    �$�Im�ےI$�pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �t   ����   �     p   ����  p    �   ?���   pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �t   ����   �     p   ����  p    �   ?���   pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �vI$�F�m��I$\     t�I$���m�$�Hp    �$�Im�ےI$�pp  �����        p           p    �           p����     ����     �������������    ?�������������   �����   "     �           �                �t  �����   �     p   ����  p    �   ?���   pp     |         p           p    �           p����  |  ����     �������������    ?�������������   �����   "     �           �                �t   �����   �     p   ����  p    �   ?���   pp    �         p           p    �           p���� �  ����     �������������    ?�������������   ��|��   "     �           �                �vI$�������I$\     t�I$���m�$�Hp    �$�Im�ےI$�pp     �        p           p    �           p����  � ����     �������������    ?�������������   ����   "     �           �                �t   �����   �     p   ����  p    �   ?���   pp     @        p           p    �           p����  @ ����     �������������    ?�������������   �����   "     �           �                �t   �����   �     p   ����  p    �   ?���   pp     @        p           p    �           p����  @ ����     �������������    ?�������������   �����   "     �           �                �q��l�����m�ۜ     t�I$���m�$�Hp    ��m��I$m��npp    8         p           p    �           p���� 8  ����     �������������    ?�������������   �����   "     �           �                �s�����������     p   ����  p    �����   ����pp    l         p           p    �           p���� l  ����     �������������    ?�������������   �����   "     �           �                �s�����������     p   ����  p    �����   ����pp    D         p           p    �           p���� D  ����     �������������    ?�������������   �����   "     �           �                �q��l�����m�ۜ     t�I$���m�$�Hp    ��m��I$m��npp    L         p           p    �           p����  l  ����     �������������    ?�������������   �����   "     �           �                �s�����������     p   ����  p    �����   ����pp    8         p           p    �           p����  8  ����     �������������    ?�������������   �����   "     �           �                �s�����������     p   ����  p    �����   ����pp     @        p           p    �           p����   @ ����     �������������    ?�������������   �����   "     �           �                �q��l�����m�ۜ     t�I$���m�$�Hp    ��m��I$m��npp      @        p           p    �           p����  @ ����     �������������    ?�������������   �����   "     �           �                �s�����������     p   ����  p    �����   ����pp      �        p           p    �           p����  � ����     �������������    ?�������������   ����   "     �           �                �s�����������     p   ����  p    �����   ����pp              p           p    �           p���� �  ����     �������������    ?�������������   �����   "     �           �                �q��l�����m�ۜ     t�I$���m�$�Hp    ��m��I$m��npp     <         p           p    �           p����  @  ����     �������������    ?�������������   �����   "     �           �                �s�����������     p   ����  p    �����   ����pp               p           p    �           p����     ����     �������������    ?�������������   �����   "     �           �                �s�����������     p   ����  p    �����   ����pp               p           p    �           p����    ����     �������������    ?�������������           "     �           �                �q��l    m�ۜ     t�I$���m�$�Hp    ��m��I$m��npp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �s����   ?���     p   ����  p    �����   ����pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �s����   ?���     p   ����  p    �����   ����pp                p           p    �           p�������������     �������������    ?�������������           "     �           �                �q��m�$�Im�ۜ     t�I$���m�$�Hp    ��m��I$m��npp                p           p    �           p�������������     �������������    ?�������������������������     �           �    ?������������p                p   ����  p    �           p������������     p           p    ��������������                �������������                �                �           �                ������������     p   ����  p    �������������������������     p           p    ��������������                �������������                �                �           �                ������������     t�I$���m�$�Hp    �������������������������     p           p    ��������������                �������������                �                �           �                ������������     p   ����  p    �������������������������     p           p    ��������������                �������������                �                �           �                ������������     p   ����  p    �������������                  p           p                  �������������     �������������    ��������������������������     �           �    �������������                  sm��rI$�6�m�p                                    p           p                  �������������     �������������    ��������������������������     �           �    �������������                  w����   ���p                                    p           p                  �������������     �������������    ��������������������������     �           �    �������������                  w����   ���p                                    p           p                  �������������     �������������    ��������������������������     �           �    �������������                  sm��rI$�6�m�p                                    p           p                  �������������     �������������    ��������������������������     �           �    �������������                  w����   ���p                                    p     �     p                  �������������     ������������    ��������������������������     �     �     �    �������������                  w���� � ���p                                    p    d     p                  �������������     �������������    ��������������������������     �    �     �    �������������                  sm��rK��6�m�p                                    p    �     p                  �������������     ������������    ��������������������������     �    �     �    �������������                  w����� ���p                                    p    �     p                  �������������     �������������    ��������������������������     �         �    �������������                  w����� ���p                                    p    �    p                  �������������     �����������    ��������������������������     �    ��    �    �������������                  sm��rO��6�m�p                                    p    ��    p                  �������������     ������������    ��������������������������     �    �    �    �������������                  w���������p                                    p    ��    p                  �������������     ������������    ��������������������������     �    �    �    �������������                  w���������p                    ?��������       p    �    p       ���������  ���       ��     ������������    ��        �����       ��     �    �    �    ��        ��  ?��������       sm��rO'�6�m�p       ���������    ?��������       p    �    p       ���������  ���       ��     ������������    ��        �����       ��     �    �    �    ��        ��  ?��������       w��������p       ���������    ?��������       p         p       ���������  ���       ��     �������������    ��        �����       ��     �         �    ��        ��  ?��������       w���� ���p       ���������    ?��������       p    �     p       ���������  ���       ��     �������������    ��        �����       ��     �         �    ��        ��  ?��������       sm��rO��6�m�p       ���������    ?��������       p     �     p       ���������  ���       ��     ������������    ��        �����       ��     �    �     �    ��        ��  ?��������       w����� ���p       ���������    ?��������       p     p     p       ���������  ���       ��     ������������    ��        �����       ��     �     �     �    ��        ��  ?��������       w���� � ���p       ���������    ?��������       p           p       ���������  ���       ��     �������������    ��        �����       ��     �           �    ��        ��  ?��������       sm��rI$�6�m�p       ���������    ?��������       p           p       ���������  ���       ��     �������������    ��        �����       ��     �           �    ��        ��  ?��������       w����   ���p       ���������    ?��������       p           p       ���������  ���       ��     �������������    ��        �����       ��     �           �    ��        ��  ?��������       w����   ���p       ���������    ?��������       p           p       ���������    @              �������������                  @              �           �                  ?��������       sm��rI$�6�m�p       ���������    ?��������       p           p       ���������    @              �������������                  @              �           �                  ?��������       w����   ���p       ���������    ?��������       p           p       ���������    @              �������������                  @              �           �                  ?��������       w����   ���p       ���������    ?��������       p           p       ���������    @              �������������                  @              �           �                  ?��������       sm��rI$�6�m�p       ���������    ?��������       p           p       ���������    @              �������������                  @              �           �                  ?��������       w����   ���p       ���������    ?��������       p           p       ���������    @              �������������                  @              �           �                  ?��������       w����   ���p       ���������    ?��������       p           p       ���������    @              �������������                  @              �������������                  ?��������       p           p       ���������    ?��������       ������������       ���������    @              �                             @              �                             ?��������       ������������       ���������    ?��������       ������������       ���������    @              �                             @              �                             ?��������       ������������       ���������                    ������������                    ��������       �                 ���������    ��������       �                 ���������                    ������������                                                                     ��������       �������������      ���������    ��������       �������������      ���������                                                                                                      ��������       �������������      ���������    ��������       �������������      ���������                                                                                                      ��������       �������������      ���������    ��������       �������������      ���������                                                                                                      ��������       �������������      ���������    ��������       �������������      ���������                                                                                                      ��������       �������������      ���������    ��������       �������������      ���������                                                                                                      ��������       �������������      ���������    ��������       �������������      ���������                                                                                                      ��������       �������������      ���������    ��������       �������������      ���������                                                                                                      ��������       �������������      ���������    ��������       �������������      ���������                                                                                                                                                       