��a  �8�G                    |�      �0 �                                     |�      �0 �                                     |�      �0 �                                     |�      �0 �                                     ��         �                                     ��         �                                     ��         �                                     ��         �                                     ��         �                                     ��         �                                     ��         �                                     ��         �                                     ������y�7�y��                                    ������y�7�y��                                    ������y�7�y��                                    ������y�7�y��                                    ��6ـ7`�7l�0                                    ��6ـ7`�7l�0                                    ��6ـ7`�7l�0                                    ��6ـ7`�7l�0                                    �͛3��`}�6l}��                                    �͛3��`}�6l}��                                    �͛3��`}�6l}��                                    �͛3��`}�6l}��                                                                                                                                          �͛1�6`Ͱ6l��                                                                                                                                                                                              �͛6ك6`Ͱ6lͳ0                                                                                                                                                                                             |����`}�6f}���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �                                                 �                                                 |                                                  8                                     ?�          ��                                    @           ��                                    �          �                                                  �                                   ��          }�                                             �        >                          �          ��                                              �        -�             �          ��          ��                                              8�        ?�             �          �x          ��                                                8�        88                       ��          ��        �            ��           ?�          �p        88                      _8          ��                                               �`        ;�           ��          ��          ��        �           ��          �          ��        7�           ��          ?�          �p        �           ��           ?�          �0        98           �           ��          5�X        0           �            ��          1�        n�           ���          �          ��                    �            �          �        �           ���          ��          ��        P           ���          	��          ��        ��           ���          ��          ;Ǹ                   ���           ��          ��       ��            ���         ��          ?��       �/            ���         ��          7��        7�           ���          )�          	�                      ���           )�          �        ��            ���         ��          ?��       p            ���                    $�H        ��           ��          ��          )�                     ��                        |        �v           ���          ��          ��       ��           ���                     '�        li              t�         ��          �0                        0                        |        �            ��Ӏ         2�          ��       G�           ����         �          7��        �              }          2�                                                            8        �            ��          �$          ��       ��           � �          ��          ;��        x9            �|�                     @                                                           @D           � "          @L          '��        ��              7          ��          ��        p           ���                     $ H         @                                                 c�            0           �          ��        S�            )�          ��          �p        /�            �                      �        �                                                 0                       �8          �P                     ��           �          |�        7�                                 �                                                                                      �p          }�        �             �           ?�          ��                                   �0          |                                                                                        �          �@                                    �           ��                                    `�           @                                                                                                  }�                                     �           �                                                �                                                                                                    �                                                                                                     �                                                                                                     8                                                                                                     8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 � � `     �   �    `�   �         >  � �                                                                                                                                                         � �   ` �    0 � `�   0 �  x     3  � `                                                                                                                                                         f �   `  �  �  0 � ` �   0 �       3  �  `                                                                                                                                                         f<�nlsǛ �  ��<y��9�l �   7<y�p     3sǝ�� `                                                                                                                                                         ffٳll`l� �  ��fͱ�m��x�   �f��`     >f`��6 �                                                                                                                                                         <~ٰllc� �   ��f���1��p    6~}��`     3g�ٛ��                                                                                                                                                         <`ٰllfl �   �f�����x    6`͙�`     3fٛ                                                                                                                                                          fٳl8fl� �   a�fͰ�m��l    6f͙�`     3flٛ6                                                                                                                                                          <�f03癀�   `�<y��8Ϟf�   �<|ٞ`     >c�͙��                                                                                                                                                              0              �                                                                                                                                                                                            �             �                                                                                 