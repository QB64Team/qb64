� h  X  ��������������������������p��p��p��p��0��0��0��0������������������0��0��0��0� p� p� p� p� �� �� �� ������������������������������������������?��?��?��?��������������������������������������������������������������������� �     �    �    �    �    �    �                            � � � � � � � � @ ` �   .� .�     ]  ]� >@   �  �  |� 8 t v  �  p � � �  � � � � � � � � � @ ` �   .� .�     ]  ]� >@   :  ;  |� 8  4  6  9  0                                              �    ?� �    ?� }�   ?� 8    ?�v    ?�