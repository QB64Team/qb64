��d   �qJ                                                                              ��������������                               ��������������                                                                              �������������                                              �                                            �                                �������������                         ?�      �������������                        @                    �                        ?�                   �                       @       �������������                         ?�      �������������                        @
                    �                        ;�                   �                       @       �������������                     �  ?�      �������������                       a`                   �                    �  ?�                   �                      a`      �������������                     �  ?�                                        �a `      ��������������                    �  ?�      ��������������                     �a `                                       �  �                                        �� `      ��������������                    �  �      ��������������                     �� `                                       �                                          ���      ��������������                    �        ��������������                     ���                                       �                                          �� �      ��������������                    �         ��������������                    A�� �                                       �   �                                      "��@�      ��������������                    <   �     ��������������                    #���@�                                       ?�=x�                                       ��     ��������������                    ><=x�     �           �                    �����     x   ����  �                     �}p�                                       ႏ�     ��������������                    �}p�     �           �                     ����     x   ����  �                     ���                                      �O�`     ��������������                    � ��     �           �                    ����`     #m��rI$�6�m�'                     �  �                                      8�O��     ��������������                    �   �     �           �                    8�O��     ����   ���                     �  �                                      |�G�H     ��������������                    �   �     �           �                    |�G�x     ����   ���                        �                                     ~��G� �    ��������������                       �     �           �                   ��G�0�    #m��rI$�6�m�'                      >  w�                                     ~������    ��������������                     >  �     �           �                   ���È�    ����   ���                       >  ��                                     ~qɜ��      ��������������                      6  �     �           �                   ~q���      ����   ���                       >  ��                                     �����      ��������������                      >  �     �           �                   ����      #m��rI$�6�m�'                         ��           �                         ���      �������������                        8�     �     �     �                   �㉛8     ���� � ���                      �  p          d                         �����     ��������������                             �    �     �                   ��ӑ�     ����� ���                     �             �                          ����p     �������������                              �    �     �                    ���     #m��rO��6�m�'                     �   �         �                          �����     ��������������                     @   �    �         �                   �G����    ����� ���                    ?�   q�         �                         ��� ��     ������������                   ?  �   q�    �    ��    �                    q��� ���    ���������                    >�   ��         ��                         ���'�      �������������                   >  @   ��    �    �    �                   0`�G�'� �    #m��rO��6�m�'                    x�  �          ��                         ����S�    �������������                   x    �     �    �    �                   xd���S�    ���������                      �  �          �                        �w���     �������������                         �     �    �    �                   �h�� 8    ��������                    �    �8         �                        �=���S     �������������                   �     �8    �    �    �                   ��?���S8    #m��rO'�6�m�'                   �   � �                                  ������    ��������������                  �      �    �         �                  �����|�    ���� ���                   �   � p         �                         �������    ��������������                  �      p    �         �                  �����<��    ����� ���                   �  ��            �                         ;����w��    �������������                  �  �       �    �     �                  ����9w��    #m��rK��6�m�'                   �  ��           p                         ?�����     �������������                  �  �      �     �     �                  ���� 0�    ���� � ���                     8� �                                    �����     ��������������                    (�  �    �           �                  ��� `�    ����   ���                     |�                                     ��ҟ���     ��������������                     �      �           �                  �ҟ���    #m��rI$�6�m�'                     �� >                                      �}�����    ��������������                    ��       �           �                   ������    ����   ���                    ��  �                                    �������    ��������������                   �  �   �           �                   �����ǀ   ����   ���                      ��  �                                  �������    ��������������                     (�  �   �           �                  ��9����   #m��rI$�6�m�'                     �    �                                  0�}ܿ���    ��������������                    �    �   �           �                  >�ܿ����   ����   ���                     |   > �                                   ��������    ��������������                          �   �           �                  .���������   ����   ���                     8   �                                  @l������    ��������������                    (     �   �           �                  N|�������   #m��rI$�6�m�'                       �� �                                  |�ȟ��@   ��������������                       #� �   �           �                  |�Ȝ\��   ����   ���                      w� �                                   ��G���@   ��������������                      w� �   �           �                   ��F����   ����   ���                   �   /� �                                   ��y��p@   ��������������                  �   /� �   �           �                   ��y��s�   \�I$���m�$�H�                      � �                                  ����� @   ��������������                      � �   �           �                  ������   x   ����  �                   >  >  ?� �                                  0���/�  `   ��������������                       ?� �   �           �                  >���/�  �   x   ����  �                   ?    ?� �                                  0������ `   ��������������                       >> �   �           �                  ?��������   \�I$���m�$�H�                   ?   ?� `                                  8���?� `   ��������������                      >> �   �           �                  ?���?���   x   ����  �                   ? 8�?� `                                  8�����  `   ��������������                   8   >> �   �           �                  ?ǔ����   x   ����  �                   ? |>��� `                                  8�����!� `   ��������������                   |  ?� �   �           �                  ?���rB!��   \�I$���m�$�H�                   ?�|��� `                                  <������ `   ��������������                  �|  � �   �           �                  ?����R ��   x   ����  �                   ?�|  �� `                                  <���� `   ��������������                  �|  � �   �           �                  ?����@�   x   ����  �                   ?�8   � `                                  >C���� `   ��������������                  �8   � �   �           �                  ?�C�����   \�I$���m�$�H�                   ?�    � `                                  > ����� `   ��������������                  �    � �   �           �                  ?�������   x   ����  �                   ?�       8`                                  ?���?�  `   ��������������                   �       ?�   �           �                  ?����?� ?�   x   ����  �                   ?�       8�                                  ??��?�  �   ��������������                   �       ?    �           �                  ?�?��?� ?�   \�I$���m�$�H�                   ?�      ��                                  ?� }܂�  �   ��������������                   x       �    �           �                  ?� }܂� ��   x   ����  �                   ?�       ��                                  ?� a��� �   ��������������                   8       �    �           �                  ?� a�����   x   ����  �                   �  8   ��                                  � A���� �   ��������������                   <  8   �    �           �                  � A������   \�I$���m�$�H�                   �  |   ��                                  � ��?���   ��������������                     |   �    �           �                  � �������   x   ����  �                   �� �   �                                  �  �|�@�   ��������������                   � �   �    �           �                  �� �|�O��   x   ����  �                   �� �   �                                  � �p� �   ��������������                   � �   �    �           �                  ���p���   \�I$���m�$�H�                   �� �   >�                                  �  `� �   ��������������                   � �   ?�    �           �                  �� `�?��   x   ����  �                   �� |   |�                                  �  @� �   ��������������                   � |   �    �           �                  �� @���   x   ����  �                   �| 8  ��                                  � �� �   ��������������                   � 8  ��    �           �                  �������   \�I$���m�$�H�                   �    �                                   �   �     ��������������                    �    ��    �           �                  ��  ���    x   ����  �                   ���   �                                   ��  ��     ��������������                    �   ��    �           �                  ��� ����    x   ����  �                   ���   ?                                    ��  �      ��������������                    �   ?��    �           �                  ��� �?��    \�I$���m�$�H�                   ��  �                                    ��          ��������������                    ?�  ���    �           �                  ���  ���    x   ����  �                   ��  �p                                   ��     p    ��������������                    �  ���    �           �                  ���  ���    x   ����  �                   ��� ���>                                   ��    �>    ��������������                    �� ��?�    �           �                  ���� ����    \�I$���m�$�H�                   ������<                                   ��   �<    ��������������                    �����    �           �                  ���������    x   ����  �                   ������< |                                   ���   < |    ��������������                    ������    �           �                  ���������    x   ����  �                    ��  � �                                    ��  � �    ��������������                    �����     �           �                   ���������    #m��rI$�6�m�'                    �� ��                                    �� ��    ��������������                    ���?�     �           �                   ��������    ����   ���                    � ��� �                                    � ��� �    ��������������                    �  ��     �           �                   ��������    ����   ���                    ?� �� �                                    ?� �� �    ��������������                     �� ��     �           �                   ?��������    #m��rI$�6�m�'                    ��    �                                    ��    �    ��������������                     �����     �           �                   ��������    ����   ���                    ��    ?�                                    ��    ?�    ��������������                     �����     �           �                   ��������    ����   ���                    ��    �                                    ��    �    ��������������                     �����     �           �                   ��������    #m��rI$�6�m�'                    ��   �                                     ��   �     ��������������                     ����      �           �                   �������     ����   ���                      ~                            ����������������   ����������������������     ����������������������������           �                     ���       ����   ���      ����������������  �������                                  ��  �       ��������������                     �?���       �           �     �������������������������#m��rI$�6�m�'      ?����������������  �������                  @               ��  �       ��������������     @               ����       �           �     ?�����������������������������   ���      ������������������������                  �               ����       ��������������     �               � ��       �           �     �����������������������������   ���      ��������������������������                                 �����       ��������������                    �   �       �           �     ��������������������������#m��rI$�6�m�'     �              ���p                        �����������������������������������������    ����������������   ���������           �    �              ���p       ����   ���     �              ���p                        �����������������������������������������    ����������������   ���������           �    �              ���p       ����   ���     �              ���p                        '�����������������������������������������    '����������������   ���������           �    �              ���p       #m��rI$�6�m�'     �              ?���p                        G�����������������������������������������    G����������������   ���������           �    �              ?���p       ����   ���     x              ���p                         ������������������������������������������     ������������������ ���������           �    x              ���p       ����   ���     >�              ���p                        A�����������������������������������������    A              �� �                   �    >��rI$�6�m�$�I#m����r6�m�$�I#m��rI$�6�m�'     }�               G��p                        �����������������������������������������    �              �x8 �                   �    }���   ���   �� ��p���   ����   ���     ��               �� p                       ?����������������> ����������������������                  ��� �                   �    ����   ���   �� �� p���   ����   ���    ��               �� p                       �����������������~ ����������������������   @              �_� �                   �   ���rI$�6�m�$�I#m� �� r6�m�$�I#m��rI$�6�m�'    �                �� p                       ������������������� ����������������������   �              �? �                   �   ���   ���   ���� p���   ����   ���    �               �� p                       !�����������������? ����������������������   !               ��� �                   �   ����   ���   ���� p���   ����   ���    �               �� p                       C�����������������������������������������   B               ����                   �   ���rI$�6�m�$�I#m����r6�m�$�I#m��rI$�6�m�'    x               ���p                        ������������������`�����������������������    �               �����                   �   {���   ���   �����p���   ����   ���    >�               ���p                       A������������������������������������������   A               �x? �                   �   >����   ���   �����p���   ����   ���    }�               ��p                       �����������������������������������������   �               ��ƀ�                   �   }��rI$�6�m�$�I#m����r6�m�$�I#m��rI$�6�m�'    ��               ߎ�p                      ?�����������������@�����������������������                  ��� �                   �   �����   ���   �����p���   ����   ���   ��               ��p                      ������������������������������������������  @               �x?��                   �  �����   ���   �����p���   ����   ���   �                ~��p                      ������������������8�����������������������  �               ��ƀ�                   �  �I$���m�$�H�m�ܒG~���u�$�H�m�ܒI$���m�$�H�   �                }ߎ�p                      !������������������@�����������������������  !                ��� �                   �  �   ����  ���� }���w�  ����   ����  �   �                ��p                      C�������������������������������������������  B                �x?��                   �  �   ����  ���� ���w�  ����   ����  �   x                ~��p                       �������������������8�����������������������   �                ��ƀ�                   �  x�I$���m�$�H�m�ܒG~���u�$�H�m�ܒI$���m�$�H�   >�                }ߎ�p                      A������������������@�����������������������  A                ��� �                   �  >�   ����  ���� }���w�  ����   ����  �   }�                �p                      ��������������������������������������������  �                ����                   �  }�   ����  ���� ��w�  ����   ����  �   ��                ~��p                     ?������������������0�����������������������                  ����                   �  �ܒI$���m�$�H�m�ܒG~���u�$�H�m�ܒI$���m�$�H�  ��                }?��p                     ������������������������������������������ @                �� �                   � ��   ����  ���� }?��w�  ����   ����  �  �                 ~��p                     ������������������� ����������������������� �                � ��                   � �x   ����  ���� ~���w�  ����   ����  �  �                 }�p                     !������������������������������������������� !                 ����                   � �ܒI$���m�$�H�m�ܒG}�u�$�H�m�ܒI$���m�$�H�  �                 {��p                     C�������������������?�@���������������������� B                 �?�@�                   � ��   ����  ���� {��w�  ����   ����  �  x                 { �p                      ���������������������@����������������������  �                 ��@�                   � {�   ����  ���� { �w�  ����   ����  �  >�                 v  �p                     A�������������������� ���������������������� A                 �� �                   � >�ܒI$���m�$�H�m�ܒGv  �u�$�H�m�ܒI$���m�$�H�  }�                   @p                     �������������������������������������������� �                 ����                   � }��   ����  ����   @w�  ����   ����  �  ��                 �  ?�                    ?������������������ ����������������������                   �                   � ���   ����  ���� �  ?��  ����   ����  � ��                 �  ?�                    ������������������  ����������������������@                   �                   ���ܒI$���m�$�H�m�ܒG�  ?��$�H�m�ܒI$���m�$�H� �                  �  �                    �������������������  �����������������������                   �                   ���   ����  ���� �  ��  ����   ����  � �                  �  �                    !�������������������  `���������������������!                    `                   ����   ����  ���� �  ��  ����   ����  � �                                            C��������������������  ����������������������B                  �  �                   ���ܒI$���m�$�H�m�ܒ@    �$�H�m�ܒI$���m�$�H� x                                             ���������������������  ���������������������� �                  �  �                   �{��   ����  ����      �  ����   ����  � >�                                            A��������������������������������������������A                  �  �                   �>���   ����  ����   � �  ����   ����  � }�                   ���                     �����������������������������������������������                  �  �                   �}�ܒI$���m�$�H�m�ܒ@����$�H�m�ܒI$���m�$�H� {�                                            �?����������������������������������������������                   �  �                   �{���   ����  ����   ���  ����   ����  � w�                                            �����������������������������������������������@                                           �w���   ����  ����   ����  ����   ����  � w                                             �������������������������������������������������                                           �wm�ܒI$���m�$�H�m�ܒI$���m�$�H�m�ܒI$���m�$�H� v                                             ������������������������������������������������                                            �v���   ����  ����   ����  ����   ����  � t                                             ������������������������������������������������                                            �u���   ����  ����   ����  ����   ����  � p                                             ������������������������������������������������                                            �sm�ܒI$���m�$�H�m�ܒI$���m�$�H�m�ܒI$���m�$�H� p                                             ������������������������������������������������                                            �w���   ����  ����   ����  ����   ����  � p                                             ������������������������������������������������                                            �w���   ����  ����   ����  ����   ����  � p                                             ������������������������������������������������                                            �t�I#m��rI$�6�m�$�I#m��rI$�6�m�$�I#m��rI$�6�m�' p                                             ������������������������������������������������                                            �p  ����   ���   ����   ���   ����   ��� p                                             ������������������������������������������������                                            �p  ����   ���   ����   ���   ����   ��� p                                             ������������������������������������������������                                            �t�I#m��rI$�6�m�$�I#m��rI$�6�m�$�I#m��rI$�6�m�' p                                             ������������������������������������������������                                            �p  ����   ���   ����   ���   ����   ��� p                                             ������������������������������������������������                                            �p  ����   ���   ����   ���   ����   ��� p                                             ������������������������������������������������                                            �t�I#m��rI$�6�m�$�I#m��rI$�6�m�$�I#m��rI$�6�m�' p                                             ������������������������������������������������                                            �p  ����   ���   ����   ���   ����   ��� p                                             ������������������������������������������������                                            �p  ����   ���   ����   ���   ����   ��� p                                             ������������������������������������������������                                            �t�I#m��rI$�6�m�$�I#m��rI$�6�m�$�I#m��rI$�6�m�' p                                             ������������������������������������������������                     �                     �p  ����   ���   ����   ���   ����   ��� p                     �                      �����������������������������������������������                     0                     �p  ����   ���   �����  ���   ����   ��� p                     ?�                      �����������������������������������������������                     �                     �t�I#m��rI$�6�m�$�I#m��?�$�6�m�$�I#m��rI$�6�m�' p                     ��                      ���������������������� ������������������������                                          �p  ����   ���   �����  ���   ����   ��� p                    ��                      ����������������������  ������������������������                      �                    �p  ����   ���   �����  ���   ����   ��� p                    ��                     ����������������������������������������������                    �@                     �t�I#m��rI$�6�m�$�I#m�����6�m�$�I#m��rI$�6�m� p                    ��                    > ����������������������?������������������������                    ?�@                    A�p  ����   ���   ����� ���   ����   ���> p                     �                    } ������������������������?�����������������������                    ��                     ��p  ����   ���   ��� � ���   ����   ���} p                     �                    � ����������������������������������������������                   ����                  �t�I#m��rI$�6�m�$�I#m���6�m�$�I#m��rI$�6�m�� p                   ��                  � ���������������������������������������������                   ���                  �p  ����   ���   ��������   ����   ���� p                   �?�                  � ���������������������������������������������                   ���                  �p  ����   ���   ����?����   ����   ���� p                   �?�                  � ��������������������� ��������������������� ��                   ���                   �t�I#m��rI$�6�m�$�I#m����?�6�m�$�I#m��rI$�6�m�� p                   � p                  � ���������������������� ����������������������@��                   �����                  @�p  ����   ���   ���� p���   ����   ��� p                   �� p                   �����������������������������������������������                   ����                   ��p  ����   ���   ���� p���   ����   ��� p                   � p                  >� ����������������������0���������������������� ��                   �����                  A �t�I#m��rI$�6�m�$�I#m����r6�m�$�I#m��rI$�6�m�� p                   � p                  }� ����������������������@���������������������� ��                   �����                  � �p  ����   ���   �����p���   ����   ��}� p                   �> p                  �� �������������������������������������������� ��                   ����                  �p  ����   ���   �����p���   ����   ���� p                   �? p                 �� ���������������������� ��������������������� ��                   �����                  �t�I#m��rI$�6�m�$�I#m����r6�m�$�I#m��rI$�6�m�� p                   ��p                 �� ���������������������� ��������������������� ��                   ����                  �p  ����   ���   �����p���   ����   ���� p                   ���p                 �� �������������������������������������������  ��                   ���                   �p  ����   ���   �����p���   ����   ���� p                   �~@p                 �� ����������������������0���������������������@ ��                   ��翈                 @ �sm�ܒI$���m�$�H�m�ܒG���u�$�H�m�ܒI$���m�$��� p                   �?@p                 � ����������������������@���������������������� ��                   �����                  � �w���   ����  ���� ���w�  ����   ���� � p                   �@p                 >�� ��������������������������������������������  ��                   ����                 A  �w���   ����  ���� ���w�  ����   ���� >�� p                   �@p                 }�� ���������������������� ���������������������  ��                   �����                 �  �sm�ܒI$���m�$�H�m�ܒG���u�$�H�m�ܒI$���m�$}�� p                   ��p                 ��� ���������������������� ��������������������  ��                   ���?�                  �w���   ����  ���� ���w�  ����   ���� ��� p                   ���p                ��� ������������������������������������������  ��                   ��?�                  �w���   ����  ���� ���w�  ����   ������� p                   �@p                ��� ����������������������0��������������������  �                   �����                  sm�ܒI$���m�$�H�m�ܒG���u�$�H�m�ܒI$���m�#��� p                   ~��p                ��� �������������������������������������������   �                   �?� �                   w���   ����  ���� ~���w�  ����   ������� p                   y�p                ��� ���������������������� ��������������������@  �                   �����                @  w���   ����  ���� y���w�  ����   ������� p                   ��p                �� ���������������������� ���������������������  �                   ��� �                 �  sm�ܒI$���m�$�H�m�ܒG���u�$�H�m�ܒI$���m��� p                   �p                >��� ���������������������� ��������������������   �                   �����                A   w���   ����  ���� ���w�  ����   ����>��� p                   x�p                }��� �������������������������������������������    �                   �?���                �    w���   ����  ���� x���w�  ����   ����}��� p                   ��p                ���� ����������������������?�������������������  @ �                   ����                 @ sm�ܒI$���m�$�H�m�ܒG���u�$�H�m�ܒI$���m����� p                   ��p               ���  ���������������������� �������������������  � �                   ��� �                 � w���   ����  ���� ���w�  ����   �������  p                   {��p               ���  ���������������������� �������������������   �                   ��� �                  w���   ����  ���� {���w�  ����   �������  p                   }�p               ���  ���������������������� �������������������    �                   �����                   sm�ܒI$���m�$�H�m�ܒG}���u�$�H�m�ܒI$���m����  p                   ~�p               ���  ������������������������������������������@   �                   ����               @   w���   ����  ���� ~���w�  ����   �������  p                   �p               ��  ����������������������@��������������������   �                   �����                �   w���   ����  ���� ���w�  ����   ������  p                   �p               >���  ����������������������0�������������������    �                   ��瀈               A    sm�ܒI$���m�$�H�m�ܒG���u�$�H�m�ܒI$���m����  p                   ��p               }���  �����������������������������������������     �                   ����               �     w���   ����  ���� ���w�  ����   ���}���  p                   �p               ����  ���������������������� ������������������  @  �                   �����                @  w���   ����  ���� ���w�  ����   �������  p                   �p              ���   ���������������������� ������������������  �  �                   �����                �  sm�ܒI$���m�$�H�m�ܒG���u�$�H�m�ܒI$���m���   p                   {��p              ���   ���������������������� ������������������    �                   ��� �                  w���   ����  ���� {���w�  ����   ������   p                   }��p              ���   ���������������������� � ����������������     �            ����������� ����������������     w���   ����        }���p              ���   p            �������~��������������������   ��������������       � � �               @    �            �       ��� �               @    sm�ܒI$���m�$�������~���������������������   p            �������������������������   ��������������       � � �               �    �            �       �� �               �    w���   ���� ��������������������������   p            ����������������������������   ��������������       � � �                   �            �       �p �                   w���   ���� ����������������������������   p            p       ���                ���   ����������������������� ����������������      �            ���������   ����������������      sm�ܒI$���m�$p       ���                ���   p            p       ���                ���   ����������������������   ����������������  @   �            ���������   ����������������  @   w���   ���� p       ���                ���   p            p       ���                ��    ����������������������   ����������������  �   �            ���������   ����������������  �   w���   ���� p       ���                ��    p            p       ���                ��    ����������������������   ����������������     �            ���������   ����������������     t�I#m��rI$�6�p       ���                ��    p            p       ���                ��    ����������������������   ����������������     �            ���������   ����������������     p  ����   �p       ���                ��    p            p       ���                ��    ����������������������   ����������������     �            ���������   ����������������     p  ����   �p       ���                ��    p            p       ���                ��    ����������������������   ����������������     �            ���������   ����������������     t�I#m��rI$�6�p       ���                ��    p            p       ���                ��    ����������������������   ����������������     �            ���������   ����������������     p  ����   �p       ���                ��    p            p       ���                ��    ����������������������   ����������������      �            ���������   ����������������      p  ����   �p       ���                ��    p            p       ���                ��    ����������������������   ���������������� @    �            ���������   ���������������� @    t�I#m��rI$�6�p       ���                ��    p            p       ���                �     ����������������������   ���������������� �    �            ���������   ���������������� �    p  ����   �p       ���                �     p            p       ���                �     ����������������������   ����������������     �            ���������   ����������������     p  ����   �p       ���                �     p            p                           �     �����������������������������������������     �            ����������������������������     t�I#m��rI$�6�p                           �     p            p                           �     �����������������������������������������     �            ����������������������������     p  ����   �p                           �     p            p                           �     �����������������������������������������     �            ����������������������������     p  ����   �p                           �     p            p                           �     �����������������������������������������     �            ����������������������������     t�I#m��rI$�6�p                           �     p            p                          �     �����������������������������������������      �            ����������������������������      p  ����   �p                           �     p            p                          �     �����������������������������������������@     �            ����������������������������@     p  ����   �p                           �     p            p          ?�                     �����������������������������������������     �            �����������������������������     t�I#m��rI$�6�p         @                      p            p          ?�                     ����������������������������������������      �            ����������������������������      p  ����   �p         @                      p            p      �  ?�                     ��������������        a`                     �            �      �  ?�                     p  ����   �p        a`                     p            p      �  ?�                     ��������������       �a `                     �            �      �  ?�                     t�I#m��rI$�6�p       �a `                     p            p      �  �                     ��������������       �� `                     �            �      �  �                     p  ����   �p       �� `                     p            p      �                       ��������������       ���                     �            �      �                       p  ����   �p       ���                     p            p      �                        ��������������      �� �                     �            �      �                        t�I#m��rI$�6�p      A�� �                     p            p      �   �                    ��������������      "��@�                     �            �      <   �                    p  ����   �p      #���@�                     p            p      ?�=x�                    ��������������       ��                    �            �      ><=x�                    p  ����   �p      �����                    p            p      �}p�                    ��������������       ႏ�                    �            �      �}p�                    t�I#m��rI$�6�p       ����                    p            p      ���                    ��������������      �O�`                    �            �      � ��                    p  ����   �p      ����`                    p            p      �  �                    ��������������      8�O��                    �            �      �   �                    p  ����   �p      8�O��                    p            p      �  �                    ��������������      |�G�H                    �            �      �   �                    t�I#m��rI$�6�p      |�G�x                    p            p         �                    ��������������     ~��G� �                   �            �         �                    p  ����   �p     ��G�0�                   p            p       >  w�                    ��������������     ~������                   �            �       >  �                    p  ����   �p     ���È�                   p            p        >  ��                    ��������������     ~qɜ��                     �            �        6  �                    sm�ܒI$���m�$p     ~q���                     p            p        >  ��                    ��������������     �����                     �            �        >  �                    w���   ���� p     ����                     p            p          ��                    ��������������     ���                     �            �          8�                    w���   ���� p     �㉛8                    p            p       �  p                    ��������������     �����                    �            �                              sm�ܒI$���m�$p     ��ӑ�                    p            p      �                       ��������������      ����p                    �            �                               w���   ���� p      ���                    p            p      �   �                   ��������������      �����                    �            �       @   �                   w���   ���� p     �G����                   p            p     ?�   q�                   ��������������      ��� ��                    �            �     ?  �   q�                   sm�ܒI$���m�$p      q��� ���                   p            p     >�   ��                   ��������������      ���'�                     �            �     >  @   ��                   w���   ���� p     0`�G�'� �                   p            p     x�  �                    ��������������      ����S�                   �            �     x    �                    w���   ���� p     xd���S�                   p            p       �  �                    ��������������     �w���                    �            �           �                    sm�ܒI$���m�$p     �h�� 8                   p            p     �    �8                   ��������������     �=���S                    �            �     �     �8                   w���   ���� p     ��?���S8                   p            p    �   � �                   ��������������     ������                   �            �    �      �                   w���   ���� p    �����|�                   p            p    �   � p                   ��������������     �������                   �            �    �      p                   sm�ܒI$���m�$p    �����<��                   p            p    �  ��                     ��������������     ;����w��                   �            �    �  �                      w���   ���� p    ����9w��                   p            p    �  ��                    ��������������     ?�����                    �            �    �  �                     w���   ���� p    ���� 0�                   p            p      8� �                   ��������������     �����                    �            �      (�  �                   sm�ܒI$���m�$p    ��� `�                   p            p      |�                    ��������������     ��ҟ���                    �            �       �                     w���   ���� p    �ҟ���                   p            p      �� >                    ��������������      �}�����                   �            �      ��                      w���   ���� p     ������                   p            p     ��  �                  ��������������      �������                   �            �     �  �                  sm�ܒI$���m�$p     �����ǀ                  p            p       ��  �                  ��������������    �������                   �            �       (�  �                  w���   ���� p    ��9����                  p            p      �    �                  ��������������    0�}ܿ���                   �            �      �    �                  w���   ���� p    >�ܿ����                  p            p      |   > �                  ��������������     ��������                   �            �            �                  sm�ܒI$���m�$p    .���������                  p            p      8   �                  ��������������    @l������                   �            �      (     �                  w���   ���� p    N|�������                  p            p        �� �                  ��������������    |�ȟ��@                  �            �         #� �                  w���   ���� p    |�Ȝ\��                  p            p       w� �                  ��������������     ��G���@                  �            �        w� �                  sm�ܒI$���m�$p     ��F����                  p            p    �   /� �                  ��������������     ��y��p@                  �            �    �   /� �                  w���   ���� p     ��y��s�                  p            p       � �                  ��������������    ����� @                  �            �        � �                  w���   ���� p    ������                  p            p    >  >  ?� �                  ��������������    0���/�  `                  �            �         ?� �                  sm�ܒI$���m�$p    >���/�  �                  p            p    ?    ?� �                  ��������������    0������ `                  �            �         >> �                  w���   ���� p    ?��������                  p            p    ?   ?� `                  ��������������    8���?� `                  �            �        >> �                  w���   ���� p    ?���?���                  p            p    ? 8�?� `                  ��������������    8�����  `                  �            �     8   >> �                  t�I#m��rI$�6�p    ?ǔ����                  p            p    ? |>��� `                  ��������������    8�����!� `                  �            �     |  ?� �                  p  ����   �p    ?���rB!��                  p            p    ?�|��� `                  ��������������    <������ `                  �            �    �|  � �                  p  ����   �p    ?����R ��                  p            p    ?�|  �� `                  ��������������    <���� `                  �            �    �|  � �                  t�I#m��rI$�6�p    ?����@�                  p            p    ?�8   � `                  ��������������    >C���� `                  �            �    �8   � �                  p  ����   �p    ?�C�����                  p   �����   p    ?�    � `                  �����    ����    > ����� `                  �   �����   �    �    � �                  p  ������ �p    ?�������                  p     �    p    ?�       8`                  ����� � ����    ?���?�  `                  �   ��?��   �     �       ?�                  t�I#o������6�p    ?����?� ?�                  p     0    p    ?�       8�                  ����� 0 ����    ??��?�  �                  �   �����   �     �       ?                   p  ������ �p    ?�?��?� ?�                  p          p    ?�      ��                  �����   ����    ?� }܂�  �                  �   �����   �     x       �                   p  ������ �p    ?� }܂� ��                  p     @    p    ?�       ��                  ����� @ ����    ?� a��� �                  �   �����   �     8       �                   t�I#o������6�p    ?� a�����                  p     @    p    �  8   ��                  ����� @ ����    � A���� �                  �   �����   �     <  8   �                   p  ������ �p    � A������                  p     ��    p    �  |   ��                  ����� �� ����    � ��?���                  �   �|}��   �       |   �                   p  ������ �p    � �������                  p     ��    p    �� �   �                  ����� �� ����    �  �|�@�                  �   �x=��   �     � �   �                   t�I#o������6�p    �� �|�O��                  p     �B    p    �� �   �                  ����� �B ����    � �p� �                  �   �x=��   �     � �   �                   p  ����� �p    ���p���                  p     ��    p    �� �   >�                  ����� � ����    �  `� �                  �   ��=��   �     � �   ?�                   p  ������ �p    �� `�?��                  p     ��    p    �� |   |�                  ����� � ����    �  @� �                  �   ��}��   �     � |   �                   t�I#o������6�p    �� @���                  p     @    p    �| 8  ��                  �����   ����    � �� �                  �   �����   �     � 8  ��                   p  ������ �p    �������                  p          p    �    �                   ����� @ ����    �   �                    �   �����   �      �    ��                   p  ������ �p    ��  ���                   p          p    ���   �                   �����   ����    ��  ��                    �   �����   �      �   ��                   t�I#o������6�p    ��� ����                   p      0    p    ���   ?                    �����   ����    ��  �                     �   �����   �      �   ?��                   p  ������ �p    ��� �?��                   p     �    p    ��  �                    �����   ����    ��                         �   �����   �      ?�  ���                   p  ������ �p    ���  ���                   p           p    ��  �p                   �����    ����    ��     p                   �   �����   �      �  ���                   t�I#o������6�p    ���  ���                   p           p    ��� ���>                   �����    ����    ��    �>                   �           �      �� ��?�                   p  �     �p    ���� ����                   p            p    ������<                   ��������������    ��   �<                   �            �      �����                   p  ����   �p    ���������                   p            p    ������< |                   ��������������    ���   < |                   �            �      ������                   t�I#m��rI$�6�p    ���������                   p            p     ��  � �                   ��������������     ��  � �                   �            �      �����                    p  ����   �p     ���������                   p            p     �� ��                   ��������������     �� ��                   �            �      ���?�                    p  ����   �p     ��������                   p            p     � ��� �                   ��������������     � ��� �                   �            �      �  ��                    t�I#m��rI$�6�p     ��������                   p            p     ?� �� �                   ��������������     ?� �� �                   �            �       �� ��                    p  ����   �p     ?��������                   p            p     ��    �                   ��������������     ��    �                   �            �       �����                    p  ����   �p     ��������                   p            p     ��    ?�                   ��������������     ��    ?�                   �            �       �����                    sm�ܒI$���m�$p     ��������                   p            p     ��    �                   ��������������     ��    �                   �            �       �����                    w���   ���� p     ��������                   p            p     ��   �                    ��������������     ��   �                    �            �       ����                     w���   ���� p     �������                    p            p     ��   �                    ��������������     ��   �                    ��������������       ����                     p            p     �������                    �������������     ���  �                    �                 ���  �                    �                    ?���                     �������������     �������                    �������������      ��  ��                    �                  ��  ��                    �                    ��                      �������������      ������                    �������������      ?�����                    �                  ?�����                    �                     �                      �������������      ?������                                        ������                    ��������������      ������                    ��������������                                                     ������                                        �����                     ��������������      �����                     ��������������                                                     �����                                         �����                     ��������������      �����                     ��������������                                                     �����                                          �����                     ��������������       �����                     ��������������                                                      �����                                          ?����                     ��������������       ?����                     ��������������                                                      ?����                                          ���                      ��������������       ���                      ��������������                                                      ���                                            ���                      ��������������        ���                      ��������������                                                       ���                                            ��                      ��������������        ��                      ��������������                                                       ��                                                                     ��������������                                 ��������������                                                                                                                               ��������������                                 ��������������                                                                                                                               ��������������                                 ��������������                                                                                                                               ��������������                                 ��������������                                                                                                                               ��������������                                 ��������������                                                                                  ��������                                    ���        ���                                 ���        ���                                   ��������                                      ��������                                    ���        ���                                 ���        ���                                   ��������                                      ��������                                    ���        ���                                 ���        ���                                   ��������                                      ��������                                    ���        ���                                 ���        ���                                   ��������                                      ��������                                    ���        ���                                 ���        ���                                   ��������                                      ��������                                    ���        ���                                 ���        ���                                   ��������                                      ��������                                    ���        ���                                 ���        ���                                   ��������                                      ��������                                    ���        ���                                 ���        ���                                   ��������                                      ��������                                              �                                             �                                     ��������                                      ��������                                              �                                             �                                     ��������                                      ��������                                              �                                             �                                     ��������                                      ��������                                              �                                             �                                     ��������                                      ��������                                              �                                             �                                     ��������                                      ��������                                              �                                             �                                     ��������                                      ��������                                              �                                             �                                     ��������                                      ��������                                              �                                             �                                     ��������                                      ��������                                              �                                             �                                     ��������                                      ��������                                              �                                             �                                     ��������                                      ��������                                              �                                             �                                     ��������                                                                                     ���������                                     ���������                                                                                                                                   ���������                                     ���������                                                                                                                                   ���������                                     ���������                                                                                                                                   ���������                                     ���������                                                                                                                                   ���������                                     ���������                                                                                                                                   ���������                                     ���������                                                                                                                                   ���������                                     ���������                                                                                                                                   ���������                                     ���������                                                                                                                                   ���������                                     ���������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      