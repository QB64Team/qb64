��h  ��Q Q  g�����0   �    �                         �������   @ ?�                        ����d   ��� �      ?�                 n��?���    ?� D    ��                �������   c���                      ���  <���  H����	     `                 _�0  /�`  �<  0�  �  �             ��    ��  @      �  � @            ���   ��  `�       ��  � �    �       �A�  ���  ��  � P   ?�  �     �  �   ���  ��� ��  ��   �  �    �  �   /�`  �?� `  �  ��  ��    `  �   [��p  ��� $�p  ��  �  �`    p  �   ���  `���(	��  a�
 @�  �0   �  `   ���  �g��@�  �� �  �   �  �   o��  �3� �&�  �p� �  �    �  �   _� �  �� �l �  �2� �  �     �  �   �� �  ��� X �  � @  �  �     �  �  �� v  ;���@� v  ;��  @ �  ?�    v  ;�   ~  {  ; ?��0 {  ; @  �    �    {  ;    @ ;`v ���` ;pv �  � ?�  �    ;  v  � �� �
n �� �
�     ?p~  �     n    �� ��l �� ��� `   p~  �    pl  @ �   \  ��� ��� �   p|  `     \    �  � �  ��� ���  �   � �  `    � �    �  �L�  W�  泸  �   ��  0    �@�   �  ���  _�  �3�  �   ��  0    ���   �  � �  k�  ���  l     p        @   �  ���  +�  ���  ,   � �      � �   �  � �  /�  ���  ,   ��      � �   �  ���  �  ��  6   ���      � �   �  ���  �,  �!�  6   ?=�~        |   �  ?�~  �,  ?� �     >�>      >  >   �  >�>  �,  ? ~     |�ߟ      <     �  z@�/  �\  z�b�      }^�_      x     �  ��� 
�X  ��P�     z��       �    �  ��  �H     0  ����          �  ���  �@  X   8  �����           ���s����O����� ?���_�w��� �� � �� ���(�
���O��"�� ?��������� ��   �� �  X�  �@  "   ?���������          � (�
` �@ "`  ?���������          � S�` �@ �`  ?���_�w���     �    �  �ǈ  �@  	H   8  �����           �  ��  �H     0  ����           �  ��Ѐ �X  �P�     z��             �  zs��  �  z���      }\_      x O   �  >�.  �,  > .     }���      <     �  ?�~  �,  ?  ~     >���      >  >   �  ���  �,  � �     ?}�~        |   �  ���  �  �c�     ���      � �   �  ��  +�  ��  (   ���      ��   �  ���  /�  ���  ,   ��      ��   �  ���  /�  ���  h   ���      ���   �  ���  W�  ��  P   ���  8     ��   �   ��   _�   ��   X   ���  0     ��    �  �$  ��� t$  �   ���  p    p     �     ���    �   � �  `          �� @ 
 _�� @ 
 @   � �  �        @ �� $  � � � $  � `   � ~  �        @ ` �  ���` �  �  � ?  ~ �        � p   D ���p   D �  �   ? �       � �� �   ��@� �   �  ` ~  ?�          ��   @�� L   @  0 �  �          ��    �� 6        �  �          �� $   �o��  $   �l   �  �        �  ��@  �_���@  ��  �  �(    @   �  ����   P���@��   Q�  �  �p    �   @0  �d�  #�  d�  #`   ��  ��    �    `  =��   "�� �   "�   ��  ��   �     �  ��   �  �       �  ��    A       ��    ��   p         ?�  �     0       �   �x  �8    �   �   �            ��   7��  0  4 @   �  �         0   ���  ���  �  �    �  �     �   �   ��c��_��   c��`      �  �      `       ���?���    \?��     ?��              }������    ��       ���       ��     �������      ���        �         ?�      �������   @ �                          �������                                                                   Q Q  g�����0   �    �                         �������   @                           �����d   �     �                         n�������         D                        �������    �                         ��������  H �� 	      �                _�����`  � � �   ��              ��������  @ q���       8  @            ���  x���  ����    � p    �            ��   ?��    <  P   �  �              ��`  ��  p      �  �     `      /��`  ���  `  �   �  �      `  �   [��p  ��� $ cx  �    �  �     p  �   ��G�  u���( ǰ  u 
 @ ?�  �    �  p   ����  ����@��  �  G�  �    �  �   o�A�  �?� �q�  � � ��  ��    �  �   _���  ��� ���  à� �  �@     �  �   �� �  ���� ��  �� @ �  �      �  �   �� v  ;�_��@ v  ;��    �  ?�0    v  ;�  � {  ; ��� {� ; L       8     {  ;   � ;`v %���& ;pv &    ?�       ;  v   �� �
n �� l �
�     ?p~       n   �� ��l �� X ���      p~      pl   �  \ 	� � ��� 	�  ` p|       \   �� � � �� � ��� �  @ � �      � �   �` �L� ��p 泸 �  � �� �    �@�  � �@ ��� ��` �3� �  � �� �    ���  � �@ � � ��` ��� �  �   p �      @  � �� ��� _�� ��� `   � �  �    � �  @ �� � � �� ��� `   ��  �    � �  @ �� ��� /� � �� 0   ���  �    � �    �� ���  ��� �!� �   ?=�~  `      |    �  ?�~  ��� ?� � �   >�>  `    >  >    �  >�>  ��� ? ~  �   |�ߟ  `    <      �  z@�/  ��� z�b�  �   }^�_  `    x      �  ��� W�  ��P� �   z��  0     �    �  ��  �	    �   ���� p         �  ���  �  X     ����� �          ���s��߀����� ���_�w��� �� � �� ���(�
�߀��"�� ��������� ��   �� �  X�  �  "   ���������          � (�
` � "`  ���������          � S�` � �`  ���_�w���     �    �  �ǈ  �  	H    ����� �          �  ��  �	    �   ���� p          �  ��Ѐ �	  �P�    z��  p           �  zs��  ��  z���  �   }\_  p    x O    �  >�.  ��� > .  �   }���  p    <      �  ?�~  ��� ?  ~  �   >���  `    >  >    �  ���  ��� � �  �   ?}�~  `      |    �� ��� /�� �c� 0   ���  �    � �    �� �� _�� �� @   ���  �    ��  @ �� ��� �� ��� `   ��  �    ��  @ �@ ��� ��` ��� �  � ��� �    ���  � �@ ��� ��` �� �  � ��� �     ��  � �`  ��  ��p  ��  �  � ��� �     ��   � �� �$ �� t$    @ ��� �    p    ��   	�� �   	�  @ � �           �X @ 
 
� � @ 
 
�    � �           �� $  � �� L $  �    0 � ~           � �  &���& �  '    ?  ~           �   D i���3   D j      ?           �퀐   ���@��   �    ~  ?�8         ���  A��� 
�  A�   �  �p          ��A   _�� a   P   ��  ��        @  ���$   ���� �$   ��   ��  ��    �    ��  ��\@  ���\@  �@   ��  �    @@   �   �� �   B���@ ��   B�   �  �      �   B   ���  ��   P�       ?�  �     �      =��  ��         �  �            ��   '��  
  $    �  �             ���  8���   �� ��     �  �     �   �   �q��_�x  � q��` �    �  ?�      p      �������   ,�  @    ��             ��������   ��      ���       ��    ���������    ���        �         �      ���������     �                           }�������                                   �������                                    �������   @                             �������                                                                   Q Q  g�����0   �8  �                         �?���}�   @�  �                      ~�����d   �    @�                        n������       D                        ��������                            ���������  H@    	                        ^������`  �  �  B�  �     �             ���`���  B  �� !     �   @            ����/���   �0     � �� �            ��������  1��� P      8               ��G  q��  ���    8               /��  ��    8    �  �              [��   �� $@      �  �             ���0  ���( 0   
 @��  � �    0      ����  ����A �  � A  �  �     �  �   m���  ��� � A�  � $�  ?�  �     �  �   _��  �� � ��  ܀� a�  �      �  �   ��0�  �?�0�  �@ @ ��  ��     �  �   ��`v  ;���H`v  ;�   ��  ?��    v  ;�   ��{  ;/����{  ;0      �    {  ;    o��;`v �����;pv�    ?�  `     ;  v    �� �
n �����
� �    ?p~ p      n   �� ��l K��  ��� L   p~ 8     pl   ��  \ +��  ��� (    p|       \   �� � � ��@, ��� 6    � �      � �   �� �L� ��@, 泸     ��      �@�   � ��� ���X �3�  @  ��      ���   � � � 
���X ��� 
       p        @   � ��� ��0 ��� �  @ � �      � �   �  � � �� � ��� �  @ ��      � �   �� ��� � � ��    @ ��� �    � �   �` ��� �� ` �!� �  � ?=�~ �      |  � �` ?�~ ��` ?� � �  � >�> �    >  >  � �@ >�> ��` ? ~ �  � |�ߟ �    <    � �@ z@�/ ��` z�b� �  � }^�_ �    x    � �� ���_� � ��P�`   z��  �     �   @ �� �� ��  `   ���� �        @ �� ��� �� X `   ����� �         @ ���s�������` ��_�w���  � � �@ ���(�
����"�` ��������  �   �@ �� X�  �� "  ` ��������         @ ��(�
` o��"` p ��������         @ ��S�` o���` p ��_�w���     �   @ �� �ǈ �� 	H `   ����� �         @ �� �� ��  `   ���� �         @ �� ��Ѐ_� � �P�`   z��  �          @ �@ zs�� ��` z��� �  � }\_ �    x O  � �@ >�. ��` > . �  � }��� �    <    � �` ?�~ ��` ?  ~ �  � >��� �    >  >  � �` ��� �� ` � � �  � ?}�~ �      |  � �� ��� � � �c�    @ ��� �    � �   �  �� �� � �� �  @ ���      ��   � ��� ��0 ��� �  @ ��      ��   � ��� 
���X ��� 
     ���      ���   � ��� ���X ��  @  ���       ��   ��  ��  ��@,  ��      ���       ��    �� �$ ��@. t$ 6    ���      p    ��   /��    ,    � �           �� @ 
 K��  @ 
 L   � � 8          ��$  � ���	�$  � �    � ~ 8          o��� ������ �    ?  ~ p           w�@  D_���@  D@  �  ? �       @  �� �  ��@0�  @   �~  ?��       @  ���  M���  �  M�   ��  ��    �   �  ���   ߀ O   �    p�  �     @      ���$   ����  0$   �     ?�  �     0    �   ���@  ���� @  �    �  �     @   �   ��   �}�@��    �   �  �     �      ��    o��     p     �  �         `   =���  1���  �  q�      �  �      �  �   ��������  ��ƀ    ~  ?       0      ����;���    n�:       ��         8    {������x  � �� �    ���       ��    ���������   ���  @     �         �     ������{�  � �  �                        ���������                                   ���������                                }�������                                   �������                                   �������   @                            �������                                                                   Q Q  g�����0   �8  �                         �?���}�   @�  �                      ~�����d   �    @�                        n������       D                        ��������                            ���������  H@    	                        ^�������`  �      B�  �     �             ���������  B      !          @            ���������            �      �            ��������   �  P                       ��������  ��      �              /����?���   �0    ��               [�������� $@ ���       0               ����  1���(  G�� 
 @� 8    �            ����   ����A �  0� A   x                m��  ?�� �   0 $�  �  �            _��l  �� � l   � �  �      l      ����  ��� �  �  @ �  �      �  �   ���v  ;����H v  ;�    �  ?�     v  ;�   ��{  ;���� .{  ;;           {  ;    o��;`v���� X;pv�     ?�       ;  v    ����
n ��� ��
��    @?p~       n    ��@��l_�� p���`   �p~�     pl   ��@ \ ��� `����   �p|�      \ �  ���� ���@����p    � � �     � � @  �� �L� ���@�泸�    �� `     �@�    � ��� ����	��3� � @ �� p     ���    � � � S��� ��� T      p 8       @   � ��� S��� ��� T    � � 8     � �   �� � � /��  ��� ,    ��      � �   �� ��� +��  �� (    ���      � �   �� ��� ��  �!� 6    ?=�~        |   �� ?�~ �� , ?� �     >�>      >  >   �� >�> �� , ? ~     |�ߟ      <     �� z@�/ �� , z�b�     }^�_      x     �� ���
�� X ��P�     z��       �    �� �� 
�� X       ����          �� ��� 
�� X X      �����           ���s���� _���   ?��_�w��   � � �  ���(�
��� _�"�   ?�������   �   �  �� X� �� @ "    ?�������           ��(�
`�� @"`   ?�������           ��S�`� @�`�  ?��_�w��      �    �� �ǈ �� X 	H      �����           �� �� 
�� X       ����           �� ��Ѐ
�� X �P�     z��             �� zs�� �� , z���     }\_      x O   �� >�. �� , > .     }���      <     �� ?�~ �� , ?  ~     >���      >  >   �� ��� ��  � � 4    ?}�~        |   �� ��� +��  �c� (    ���      � �   �� �� /��  �� ,    ���      ��   � ��� S��� ��� T    �� 8     ��   � ��� _��� ��� X    ��� 0     ���   � ��� ������� � @ ��� p      ��   ��� ��  ���@� �� �    ��� `      ��     ����$O��@�t$P    ��� �     p  @  ��` �� ` `   �� ��        @  ��0@ 
��� 0@ 
�   �� ��        �  ���$  �����$  ��    `� ~     @     o�(� ��� �� �    p?  ~           w��  D6���� V  D7    8  ?          ���  m���@ +  n     �  ?�          ���  ���        �  �          ���   7�߀ 
   8     �  �            ����   ����  �   �     �  �     �   �   ���B  1?��� C  q@     �  �      @      ��y���}�@� ��΀ �    >  ?       8      ����1���    ~�2       ��         0    =��������   ��       ���       ��    ��������   ��`      ?��        �     ��������     ?��                          {�������x  �      �                       ���������         @                       ������{�  �     �                        ���������                                   ���������                                }�������                                   �������                                   �������   @                            �������                                                                   Q Q  g�����0   �8  �                         �?���}�   @�  �                      ~�����d   �    @�                        n������       D                        ��������                            ���������  H@    	                        ^�������`  �      B�  �     �             ���������  B      !          @            ���������            �      �            ���������       P                       ���������                            /���������                              [��������� $@  �                         �����?����(  ��  
 @�  �   �            �����o����A  �p  A    ��              m�������� �  8���  $�     p               _��g� ���� �  ���  �                   ����  �� �  }�  @  &               ���6  :���H 6  :@     �  =�       8    ��{  ;����� {  ;�    �  ~@     ;  :    o���`v����� �pv�     ?�        ;  v    ����
no��� ��
��     ?p~       n    �����l���  ���T    
p~(      pl    ��� \3���  .���2     p|       \    ���� ����@ L���     0� �      � �   ����L�
���@ X泸
      ��      �@�   ��������� ��3�� @ @��      ���   �@� �����P����    �  p�       @ �  �@�������`����    �� ��     � � �  ���� ���  ����@    �� �     � � @  �������� ���`    ��� �     � � @  ������_�� ��!�@    ?=�~ �       | @  ���?�~ ��� �?� � �    >�> `     >  >    �� >�> ��� �? ~ �    |�ߟ p     <      �� z@�/ ��� �z�b� �    }^�_ p     x      �� ������ ���P��    z�� 0      �    �� �� W��   X    ����0          �� ��� _��  X X    �����0           ���s���� ���   ��_�w��   � � �  ���(�
��� �"�   �������   �   �  �� X� �� 
 "    �������           ��(�
`�� 
"`   �������           ��S�`�� 
�`   ��_�w��      �    �� �ǈ _��  	H X    �����0           �� �� W��   X    ����0           �� ��Ѐ��� ��P��    z�� 0            �� zs�� ��� �z��� �    }\_ p     x O    ���>�. ��� �> . �    }��� `     <      ���?�~ ��� �?  ~ �    >��� `     >  >    ������_�� �� �@    ?}�~ �       | @  �������� ��c�`    ��� �     � � @  �������  ���@    ��� �     �� @  �@�������`����    ����     �� �  �`�������p����    �����     ��� �  ��������� ���� @ @���       ��   ��X �� 
���@ � �� 
�     ���       ��    ����$���@ Lt$     0���      p    ��� 7���  & 6     � �           ���@ 
o���  ;@ 
l    � �          ���  ����� �  ��     � ~0          o��D� ?���� D� 0     �  ~�           w��  D����   D`    �  ?�       @   ����  ����@ �  �      �  ?�      �  �   ����  b����   �  b�     |                ��������߀  x��         |             �����w����   �t       ��         p    ����������  ��      ���        ��    ��������}�@� ���  �     ?�         �     ���������     �                           =���������                                 ���������                               ���������                                  {�������x  �      �                       ���������         @                       ������{�  �     �                        ���������                                   ���������                                }�������                                   �������                                   �������   @                            �������                                                                   Q Q  g�����0   �8  �                         �?���}�   @�  �                      ~�����d   �    @�                        n������       D                        ��������                            ���������  H@    	                        ^�������`  �      B�  �     �             ���������  B      !          @            ���������            �      �            ���������       P                       ���������                            /���������                              [��������� $@                             �����������(        
 @�       �            �����������A        A                     m�������� �   �   $�                      _������� �   p�  �   �                �����o���  �p   @   ��               ����������H  ���        `              ���  �����  �        x              o���`c�����  cp�       � |         `    ����
h����  ��
�      p        h    �����m���  ���@     �p~�      pl    ���N ]����  n��ߠ     �p|@       \    ���� �_���@ N���P     �� ��      � �    ����L�����@ �泸�     ��P      �@�    �����G���� �3�D  @ ��8      ���    ��� �!���� ���"       p        @    �����7���� ���6     � �      � �   ���� ����  ,���     ��      � �    ���������  X��      ���      � �   ���������  X�!�      ?=�~        |    ���?�~��  8?� ��    @>�>      >  >   �� >�>���  �? ~�    @|�ߟ      <     ���z@�/��  �z�b�     @}^�_�     x     ������?��  ���P�@    @z���      �    ��@����� `�    ����        �  �� ������  X�    �������         �  ��?s�~��� ?�~�    ��_�w��    ? � ~�  ��?(�
~��� ?"~�    �������    ?   ~�  �� X� ���  " �    �������         �  ��(�
`��� "`�    �������         �  ��S�`��� �`�    ��_�w��      �  �  ��@�ǈ��� `	H�    �������         �  ��@����� `�    ����         �  �����Ѕ?��  ��P�@    @z���            ���zs����  �z���     @}\_�     x O   �� >�.���  �> .�    @}���      <     ���?�~��  8?  ~�    @>���      >  >   ������
���  X� �
      ?}�~        |   ���������  X�c�      ���      � �   ��������  ,��     ���      ��   �����'���� .���&     ��      ��   �����/���� ���l     ���      ���   �����s���� ��t  @ ���       ��   ������ ����@ ��� �     ���0       ��    �����%����@ �t%�     ���`     p     ���2 ���  2 `     �� ��       @   ����@ ����  �@ �     �� ��      �  �   ����  �����  �  ��      �        d      o��Ѐ ������  P��       ?  ~             w���p�����  <|      � �             �����k����@  �l       ��         `    ����������   ��      ���        ��    ����O���߀   ���        ?�         �     �����������    �                           �����������                               ��������}�@�       �                       ���������                                  =���������                                 ���������                               ���������                                  {�������x  �      �                       ���������         @                       ������{�  �     �                        ���������                                   ���������                                }�������                                   �������                                   �������   @                            �������                                                                   Q Q    <�       � �       @                  �đ�      ;n        �                 >�>`      �� ��      @                  �����               @                ;��f     �l�      �                 L�?�_�     3��f      � @�               �������    @       �  �              g�����`    �   �     @                  ����?�   �   �`                        ;�����h   �    �                       �������                @              =�������                               [�������   $  ?�    @                  ��`?�v�  H��� �      �                n���o��@  � �p D�  @  ��              }������`  � 8���  �  !   p B             ��!  b�� D ��� @                    ���  ��� @�  p�    >              ��  8_��   8`  � �  ?� �      8    
���  :/��  �  :0 P   �     ;  :    ���`v��� 	 �pv�@  ?�       ;  v    ���
nk�� 
@��
��    ?p~       n    +����l7��  7���t    @p~     pl    ;� \3�� �.���2   p|       \    W�� ��� (�\���    � �      � �    W�P�L�
� ( �泸
�@   ��      �@�   ��������	 ��3�  @ @���     ���   ��`� ����Bp����  �  p�       @ �  ��@����߀P`����   �� ��     � � �  ���� �_� R����` �� �� �     � � @  {�����_������@   ��� �     � � @  _�����_��!�@  ?=�~ �       | @  [��?�~ �����?� � �    >�> `     >  >    �� >�> �� �? ~ ��� |�ߟ p     <      �� z@�/ ��@�z�b� �  }^�_ p     x      �� ������H���P��    z�� 0      �    �� �� W��H  X    ����0          �� ��� _�� 	 X X	 H �����0           ���s����H	���   ��_�w��   � � �  ���(�
���H	�"�   �������   �   �  �� X� ��  " 	 H�������           ��(�
`��H"`   �������           ��S�`��H�`   ��_�w��      �    �� �ǈ _�� 	 	H X	 H �����0           �� �� _��H  X    ����0           �� ��Ѐ���H��P��    z�� 0            �� zs�� ��@�z��� �  }\_ p     x O    �� >�. �� �> . ��� }��� p     <      [��?�~ �����?  ~ �    >��� `     >  >    _�����O�� �P  ?}�~ �       | @  {����������c�`   ��� �     � � @  �����_� R ���` �� ��� �     �� @  ��@����߀P`����   ����     �� �  ��`������Bp����  �����     ��� �  ���������	 ���� @ @���       ��   W�X �� 
�� ( � �� 
 @   ���       ��    W��$�� (�\t$    ���      p    ;� 7�� �& 6   � �           +��@ 
o�� @@ 
l    � �          ���  ���� 
 �  ��     � ~p          ��� ?��  � 0     �  �           ��  D��    D`   �  ?�       @   ��  ��x  ��  A� �    �  ?�      �  �   ���  B���   ��      ~  ?              ��������   X��       ?  |             ����u���  ! 7�v B     ��         p    ��������  @ ��      ���        ��     ���������    ���        �         �      w�������   @ �                          /�������                                �������         @                         �������                                  �������                                   �������     @                             w�����@    �  �                          ~���      � @�                           /��o��      �                            �����       @                           �����      @                              ��o��       �                             ;���       @                                                          Q Q    <�       � �       @                  �đ�      ;n        �                 >�>`      �� ��      @                  �����               @                ;��f     �l�      �                 L�?�_�     3��f      � @�               �������    @       �  �              g�����`    �   �     @                  ����?�   �   �`                        ;�����h   �    �                       �������                @              =�������                               [�������   $        @                  ������v�  H�     �                        n������@  �  �  D�  @                   }��0��`  �  ��  �  !  �  B             ����o�� D �p @    ��               ���x��� @ �     � �              ��Ѐ ����  0��   �   |  �            
��C  !��   �  !� P  ?  ~             ���`p��� 	 �pp�@   �         p    ���
l_�� 
@�
�`     �p�       l    +�����m���  ����    @p~`     pl    ;�� \��� �ί���   p|        \    W�� �o�� (�����   � �      � �    W���L�g�� ( 7泸d @  ��      �@�    ������3���	 .�3�2  @ ��      ���    ���� ����B L���4   0  p        @   �������߀P \���     � �      � �   ��P� �
�� R ����
  ��  ��      � �   {��������� ����   @���      � �   _����� ��!�   @?=�~�       |   [�`?�~����`?� ��    �>�>�     >  > �  ��@>�>�� `? ~��� �|�ߟ�     <   �  ��@z@�/��@`z�b��  �}^�_�     x   �  ��@��󐂿��H`��P��    �z���      �  �  �����_��H�`    �����        @  �������� �X`	 H ������         @  ��s���H�`   ��_�w��     � @  ��(�
��H"`   �������       @  �� X� _��  " @	 H�������         @  ��(�
`_��H"`@   �������         @  ��S�`��H�``   ��_�w��      �  @  �� �ǈ�� @	H`	 H�������         @  �������H �@    �����         @  ��@��Ђ���H`�P��    �z���          �  ��@zs����@`z����  �}\_�     x O �  ��@>�.��  `> .��� �}����     <   �  [�`?�~���� `?  ~�    �>����     >  > �  _����� �� �   @?}�~�       |   {�0������ ��c��   @���      � �   �����
�� R X��
  ��  ���      ��   �������߀P X���     ��      ��   ���������B ,���   ���      ���   ������%���	 .��&  @ ���       ��   W�� �� k�� (  �� h @  ���       ��    W���$��� (��t$�   ���8     p    ;�� ��� �
� �   � �p           +��@ O�� @@ P    �� ��       @   ���  ���� 
 �  ��     �� �      �  �   ��D� ?��  D� @      �  �      D      ��0� ���   ����             0      ��p��x  � ,|  �    � �             ����g���   �h      ��         `    ���p���   p        ���        p     ���������  !  O�  B      ?�         �     ���������  @  �                           ���������                                   w�������   @                             /�������                                �������         @                         �������                                  �������                                   �������     @                             w�����@    �  �                          ~���      � @�                           /��o��      �                            �����       @                           �����      @                              ��o��       �                             ;���       @                                                          Q Q    <�       � �       @                  �đ�      ;n        �                 >�>`      �� ��      @                  �����               @                ;��f     �l�      �                 L�?�_�     3��f      � @�               �������    @       �  �              g�����`    �   �     @                  ����?�   �   �`                        ;�����h   �    �                       �������                @              =�������                               [�������   $        @                  ������v�  H�     �                        n�������@  �      D�  @                   }�������`  �       �  !      B             �������� D      @                      ���0��� @  ��      �               ����_���  �`   �  ��  �            
���0���   0  P  � �              �������� 	  0�� @     x              ����
b��� 
@ a�
�      p|        `    +��E��i��   ����    @ ?p~      ph    ;� ^?�� ����@    �p}�       \    W�N� ��� (�N���    �� ��      � �    W����L���� ( �泸� @  ��`      �@�    ������/���	 �3�   @ ��p      ���    ���� �W���B 
���X     p0        @   �������߀P ���    � �8      � �   ���� ��� R ���  �� ��      � �   {��������� (��    ���      � �   _������ (�!�   ?=�~        |   [��?�~���� X?� �      >�>      >  >   ���>�>��  P? ~ ��  |�ߟ      <     ���z@�/��@ Pz�b�    }^�_      x     ��Є�����H P��P�      z��       �    �� ����H ��    @����           �� �����  �X�	 H `�����            ���s�}���H ��}�    �_�w�      � }   ���(�
}���H �"}�    �����        }   ���X����  �"�	 H �����            ���(�
a���H �"a�    ~�����            ���S�a���H ��a�    ~�_�w�       �    �� �ǈ��  �	H�	 H `�����            �� ����H ��    @����            ��P��Ђ��H ЅP��     z��             ���zs����@ Pz���    }\_      x O   ���>�.��  X> . ��  }���      <     [��?�~���� X?  ~      >���      >  >   _������ ,� �   ?}�~        |   {��������� ,�c�    ���      � �   �����	�� R ��
  �� ���      ��   �������߀P ���    ��8     ��   ������S���B ���T   ���8     ���   ������/���	 ����  @ ���p      ��    W�� �� W�� (  ��!X @  �����      �� @   W��$o�� (�1v&p   �����     p @   ;�� ��� �� �    �� ��      �  �   +���@ ��� @�@ �     � �       "      ��P  ��� 
  �@ ��      ?� ~             ���  ���   l@       � �             ���  k���   l     ��         `    ������x  � ��  �    ���        ��    ���������   ���       ?�         �     ���������    ?�                           ���������  !      B                        ���������  @                               ���������                                   w�������   @                             /�������                                �������         @                         �������                                  �������                                   �������     @                             w�����@    �  �                          ~���      � @�                           /��o��      �                            �����       @                           �����      @                              ��o��       �                             ;���       @                                                          Q Q    <�       � �       @                  �đ�      ;n        �                 >�>`      �� ��      @                  �����               @                ;��f     �l�      �                 L�?�_�     3��f      � @�               �������    @       �  �              g�����`    �   �     @                  ����?�   �   �`                        ;�����h   �    �                       �������                @              =�������                               [�������   $        @                  ������v�  H�     �                        n�������@  �      D�  @                   }�������`  �       �  !      B             �������� D      @                      ��������� @                            ��������   �    �       �            
��������    p   P   �               ��������� 	  ��� @    p               ���p/��� 
@ �0      � �               +���������   ���     @ pp       p     ;�� E��� � 0���     px         @    W��� ���� (� F���     ?� �       � �    W��7�L��� (  �泸� @   G��       �@�    ���c���?���	 s�3�@  @  ����      ���    ���A� ß���B a��à    �  t�        @�   �������_�߀P ����@    � ��      � �@   ����� ���� R Ͽ���  �� ��`      � �    {���������� ����    ���p      � �    _�����_� �!�X   ?=�~0        |   [��?�~W���� ?� �P     >�>8      >  >   ���>�>/��  ? ~( �� |�ߟ      <     ���z@�//��@ z�b�,   }^�_      x     ��������H ��P�     z��       �    ��������H      ����           ���������  $X 	 H �����            ���s�u���H '�v     �_�w�      � t   ���(�
w���H '"v     �����        t   ���X����   " 	 H �����            ���(�
g���H !"f     �����            ���S�g���H !�f     �_�w�       �    ����ǈ���  $	H6 	 H �����            ��������H ,6     ����            ����Ы���H �P�     z��             ���zs��+��@ z���h   }\_      x O   ���>�.+��  > .l �� }���      <     [��?�~W���� ?  ~P     >���8      >  >   _�����W� � ��   ?}�~0        |   {���������� ��c��    ���p      � �    ��������� R ����  �� ���`      ��    ���G���_�߀P g���@    ����      ��@   ���3��֟���B 3��֠    �����      ����   �����������	 ����  @  ����      ����   W��H�!�� (  �~�!� @   w���       @>�!    W���&��� (� qt'     ?���       1p&    ;�� 	��� � ('�
     � �             +���p3��� @ |4      � �         0    ��������� 
  ���       ��       � �    ���p?���   p@        ���        p     ���������    O�       ?�         �     �������x  �  �   �                       ���������                                ���������                                 ���������  !      B                        ���������  @                               ���������                                   w�������   @                             /�������                                �������         @                         �������                                  �������                                   �������     @                             w�����@    �  �                          ~���      � @�                           /��o��      �                            �����       @                           �����      @                              ��o��       �                             ;���       @                                                          