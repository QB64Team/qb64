�:a  \]�g                     <�         0                                          <�         0                                          <�         0                                          <�         0                                          f� �    �0                                          f� �    �0                                          f� �    �0                                          f� �    �0                                          `� �    �0                                          `� �    �0                                          `� �    �0                                          `� �    �0                                          `y�<�x��y�`9ͳ�                                         `y�<�x��y�`9ͳ�                                         `y�<�x��y�`9ͳ�                                         `y�<�x��y�`9ͳ�                                         <ͳf��6��m��`                                         <ͳf��6��m��`                                         <ͳf��6��m��`                                         <ͳf��6��m��`                                         ��`�|��}��1���                                         ��`�|��}��1���                                         ��`�|��}��1���                                         ��`�|��}��1���                                                                                                                                                             ��`���͛���                                                                                                                                                                                                                        fͳf���6͛`m�6`                                                                                                                                                                                                                       <y�<`|��}�08�3Ͱ                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          �                                                        �                                                        �                                                        �                                                         ,                                                         ,                                                        �                                                                                          �          	�z         .                                ^�          ?�z�        .                                ?�          ��         �                                �          0@z                                           �          @          �                                �          ��         �                                }           ��        �                                            �                                �           B�          ��       �                   �           B�         �y�       ��                   �           =           ���        ��                    �                      �                                                     ?�            8                              ?�         ��        ���                  �                     ��         ?���                               +�         ?��        @                               A`          pp�        �[           �                ��         ���       ����          �      �          ��         ���        ����          �                            pp`       [            �       �                     ��       �K �          �      �          ?��         ?��       �P���          �       �          ��         ���       �����         H      ^                      �`        �K                   :           ?�                   n  P         �      ��         ��        ���       �����         �      ?�          ?��         ���       �����         @      @ �         @?��          `        n  P                  �           A��                  �                  ���         ���        ���       ?����         �      ���         ���        ���       �����                           ���         	          �            �     �          ��        �           �         ��    � �        ���        ���       ����        ���    ���         ����        ���       �����         ���    �        �                       �              8�          �        
̍            �          `   ��        ���~        ��       =����߀       ����   ���        ����        ���       ������       ����   8�           �          �       "                   @ X          !�       ~E                    ��   ����       ���߀       ���       ?������       � �   ����       �����       ���       ?������       ����   @ X@                      @                     ��   	�                     �!                     � ��  ���       �����       ���       ?������       ����  ����       �����       ���       ?������       �����  �                                              � �     �        �        
��                     #   8  ���x       �����       ���       ?������       ?�����  ����       �����       ���       ?������       ?�����    �                                               8     b        @�`        ?��                     D   �  =����       �����       ���       ?������       {����~  ����       �����       ���       ?������       �����  "   `       @                                      �  $ �        V�         ��                    H    a  ;����       �����       ����      ?������       ������� ?����       �����       ����      ?������       �����                                                 �    `�  ��        }�        ?��       *      �      �    @ �����      �����       ����      ?�������      ������� ?�����      �����       ����      ?�������      ������� @   @                                                H
�p        W��        _��             @        
�  w�����      ������      ����      �������     ������� �����      ������      ����      �������      �������                                                      �\       ��x        ?���      Uk           �_� � ������      ������      ���p      �������     ������8 �����      ������      ����      �������     ������� �                           �                          �  .�� @      	���       ��@      ���         ���   ������      ������      ����      �������     ������� �����      ������      ����      �������     ������� �    @                       @                          " �w�m�        
���       ?��       ���           ���� ������      ������      ����      �������     ������� ������      ������      ����      �������     �������                                                         	 �_o��      ���@       ���       ?���          /���� ������      ������      ����       ������     �������������      ������      ����       ?������     �������                                   @                  @ {���      ���       ���       ����        :���� ������      ������      ����       ������     �����s��������      ������      ����       ������     �������                                                    �  ����       ����       ���       ����         _���တ�������     ������      �����      ������     ������x�������     ������      �����      ������     ����� ��                                                    � ���o       ����       ���        ?���  �      k����`P�������     �������     �����       ������    ��������������     �������     �����       ?������    ����� ?�                                     @                  @ �����       ���� @     ���        ���  @      ����� �������     �������     �����       ������    �����o��������     �������     �����       ������    ����� �                                                      �����@     ����@      ?����       ���  `      ����� �������     �������     ����p       ������    �����W��������     �������     �����       ������    ����� �                              �                           �����@     �����     ���@        ?���       ������������     �������     �����        �����    �����K�������     �������     �����        ?�����    ����� ��     H                      @        @                   ����p      �����     ?���         ���      ������������     �������     �����        �����    �����I�������     �������     �����        �����    ����� �                                                          ����       ������      ����        ���        �����`?������      �������     �����        �����     �����I�?������      �������     �����        �����     ����� �                                                        ����       A�����      ?����         ?���      �_����������      ������     �����         ����     �����I�������      ������     �����         ?����     ����� �                                      @                  ?����        �����     ����         ���     @����@������      ?������     ������        ����     �����I�������      ?������     ������        ����     ���� �                                               �        ����       ?����       ?����         ���      @?�����������      ������      �����        ����     ����A�������      ������      ?�����        ����     ���� �                        @                               ����        ������      ����          ?��       ?����� �������     ������      �����         ���     ?����C� �����       ������      �����         ?���     ?���� � �     �                              @                 �����         ?����     ����          ��     ������ ������       �����     �����         ���     ?���� � ������        ?����     �����         ���     ���� �              �                                        �����@         ��       ?���@         ��      ������ ������        ����      ����         ���     ���� � ������         ���      ?����         ���     ���� �               �         @   @                         ����@         ��       ���           ?���    �����  �����         ���      ����          ���    �������  �����         ���      ����          ?���    �������  `                                     @                ����           �       ����          ��     �     �  �����         ���      ����          ���    �������  �����          ��      ����          ���    �������                �                                   0   ���           �        ���          ��@               ����          ��       ����          ���               ����          ��       ���          ���               `                       �                               ��             �       ���           ?�                ����          ��       ����          ��               ����           ��       ���           ?��                                         �          @                  �             ?        ��Ѐ          �                 ���           �       ����          ��                ���           ?�       ����          ��                `  @           @                                          �             �        ��           �                 ���           ?�        ����          ��                ��            �        ���          ��                  �           0         �                                             �        ��            ?�                 ?�            �        ���           �                 �            �        ���           ?�                 0                                    @                   |            �        ��            �                 �            �        ���           �                  |            �        ��            �                 �                        �                                            �         �             �                                �         ��            �                                �         �             �                                          �                                              4         �                                              |         ?�                                              <         �                                              @                                                                 �                                                       �                                                       �                                                                                                                                                                         �                                                         8                                                         �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �  �        �    0     >`��  0      �0         �0`0                                                                                                                                                                                   �        �    0     c`��  0      �0         � 0                                                                                                                                                                                   �             0     c`��  0       0         � 0                                                                                                                                                                                <����      <���     cg���Ǐ0      >s�       ��g>                                                                                                                                                                                3�ٛ0      ��f͛0     cl��7lٰ      �``       �6m�                                                                                                                                                                                ?>�ٛ0       �3f��0     cl�lٰ      �c�       �6f3                                                                                                                                                                                0f�ٛ0       �3f̓0     cl�lٰ      �f`       �6c3                                                                                                                                                                                3f�ٛ0      ٳf͛0     cl��6lٰ      ٳf`       �6m�                                                                                                                                                                                >����      �<���     >g���g�0      �>c�       �3g3                                                                                                                                                                                                �                                                                                                                                                                                                                                      �                                                                                                  