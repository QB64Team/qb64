�oh   ��F                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ���                                             ���                                             	D                                             ���                                             ���                                             ���                                             d�4                                             ��                                             ���                                             ���                                             QD                                             _߂                                             ���                                             ���                                             \E                                             _�                                             ���                                             ���                                             �T                                             ��                                             (��                                             ���                                             u�T                                             u�                                             �_�                                             ���                                             UTT                                             UP                                             ���                                             ���                                             ]�D                                             ]                                              ���                                             ���                                             �%T                                             �$                                             *��                                             ���                                             w�                                             v                                              ���                                             ���                                             UT                                             U                                             ���                                             ���                                             _��                                             X                                              ���                                             ���                                             � �                                             � �                                             '�>                                             ���                                             ��                                             p                                              ���                                             ���                                             a4                                             a2                                             ���                                             ���                                             ���                                             �                                              ?��                                             ���                                              �                                              �                                             ��z                                             ���                                            ���                                       �����  �����                                  �������������                                  �������������                                  �������������        �                          ���� �                                  ���}�  �~���        �                         �������������                             ?�    �����  �����        �                  @      �    �                           ?�    ���}�  �~���        �                  @     �����  �����                           ?�          �              �                  @
     �������������                          ;�    �����  �����        �                  @     �������������                      �  ?�    �������������    �  �                 a`      A@� 	  A      �0�0               �  ?�    ߾��  ���߾    �  �                 a`    ������ �����      �0�0               �  ?�    ������������    �  �                �a `      A@���  A      �0�0               �  ?�    ߾��  ���߾    �  �                �a `    �������������      �0�0               �  �          �w�         �  �                �� `    ������r�����      �p�0               �  �    �����t�����    �  �                �� `    ������v�����      �p�0               �      ������������    �                  ���     ���� �      �Q�p               �      ���}���~���    �                  ���    �������������      �Q�p               �       �������������    ��                 �� �     ��� �     ��qp               �       ���}���~���    ��                 A�� �    �������������     ��qp               �   �        �7�         �   |              "��@�    ������7������     �a p�              <   �   �����7�����       |              #���@�    ������7������    ��a p�              ?�=x�   �������������    �� �               ��     AA���  A      ��@s@              ><=x�   ߾�����߾    � �              �����   �������������     ����s@              �}p�   ������Ϗ�����    �>��               ႏ�     AC���  A      ��G�              �}p�   ߾������߾    �>��               ����   �������������     ����              ���        ���         �X��             �O�`   ������������    ����0              � ��   �����������    � X��             ����`   �������������    ����0              �  �   ������������    � ���             8�O��    ���� �    �ç�H              �   �   ���}���~���    �   �             8�O��   �������������    ��'�X              �  �   ������w������    �  ��             |�G�H    ��r �    >��#�$              �   �   ���}�t�~���    �   �             |�G�x   ������v�����    >��#�<                 �        ?��          �  ��            ~��G� �  �������������   ?a��#� |                �   �����  �����     �  �            ��G�0�  �������������   ?���#�|              >  w�     A���  A     �  ;��            ~������    A� 	  A   �p��a�D              >  �   ߾��  ���߾     �  ��            ���È�  ������ �����   ����a�D               >  ��     A���	  A        }�             ~qɜ��      A���  A    �8��C�                 6  �   ߾�� ����߾        �             ~q���    �������������    �8��C�                 >  ��   ������ ������        |�             �����        �� �        ?����G�                 >  �   ����   �����        �             ����    ������ ������   ?����G�                   ��    �             |             ���     �������   ?���č�                   8�   ���      ���                     �㉛8   �������������   ?����͜               �  p    �          p  8�            �����    �������    �������                     ���      ���        �            ��ӑ�   ����     ���    ������߀             �      �������������   � �   �             ����p       �            ~�����                      ������������   �     �             ���   �������������    ~�����             �   �    A�������  A   ��   �             �����     A�������  A    ~��цp               @   �  ߾��������߾   �     �            �G����  �������������   ~#�цq�            ?�   q�    A�Z��@  A   ��   8�             ��� ��     A����x  A    ?����~�             ?  �   q�  ߾����g�߾   � P   8�             q��� ���  �������g���   8�S��~��            >�   ��  ����[m�������   ��   |p             ���'�        �[m����       ?�����             >  @   ��  ���[m�������         |p            0`�G�'� �  ����[m�������   0~#���p            x�  �    �[lZ���   <��   �              ����S�   �[lZ���    ?��܏�)�            x    �   ���[lZ������   <     �             xd���S�  ����[lZ������   <2���)�              �  �    �[m����    �p   �            �w���    ��m����   ;����                   �   ����m�������          �            �h�� 8  �����m�������   4?���            �    �8  �����mҕ�����   p     �            �=���S       ��m׵��      �����)�            �     �8  ����m׵�����   p      �            ��?���S8  �����m׵�����   q�����)�           �   � �    A��lZ4D`  A   �   � |            ������    A��l[tDX  A   ������           �      �  ߾��l[tDg�߾   �      |           �����|�  �����l[tDg���   ����>��           �   � p    A�������  A   �   � 8            �������    A�������  A    ������           �      p  ߾��������߾   �      8           �����<��  �������������   ������           �  ��    ����     ���  �  ��              ;����w��     �������      ���;��           �  �     ���      ���  �  ��             ����9w��  ����     ���  �������           �  ��   !�       �  ��  �            ?�����   !�������   ����            �  �    ���      ���  �  �   �           ���� 0�  ����     ���  ��� �             8� �  #�������  � �� À           �����   #�������   �k����             (�  �  ���      ���  � �  À          ��� `�  �������������  ��c�0���            |�   �������������  � >�  ��           ��ҟ���      �������      �~�O���               �    ���      ?���  �  �   ��          �ҟ���  �������������  ��@�O����            �� >     A�������  A  � �  �            �}�����    A�������  A    ~>�����             ��     ߾�      o�߾  � A�   �           ������  �������������  �~ �����           ��  �   A������  A  � � ?��            �������    A������  A    |�����            �  � ߾�      ��߾  � �  �           �����ǀ �������������  �|�����             ��  � �������������     � ?��          �������     ������      ��w��?��              (�  � ���      ����     �  �          ��9���� �������������  ������            �    �  � � �       ?��          0�}ܿ���   � � �  �>�_�?��             �    � ���}��}��~���    I    �          >�ܿ���� �������������  ��_���            |   > �  � � �    >     �           ��������   � � �  ������                   � ���}��}��~���           �          .��������� �������������  �A������            8   � �������������      �  �          @l������                   �K����             (     � �������������          �          N|������� �������������  '�C����              �� �                     ��  �          |�ȟ��@                 >O�O��                #� �                      �  �          |�Ȝ\��                 >O�N.��             w� �                  �   �� �           ��G���@  >          �   ?��#��               w� �  >          �   �   ;� �           ��F����                  ?��#D��          �   /� �  �����������   �   � �           ��y��p@  >          �   ?��<�p8           �   /� �  >          �  �   � �           ��y��s�                  ?��<�p9�             � �   �       ��    �  � �          ����� @  ?������������  ��?�@�               � �  >          �   �   � �          ������  �����������   ��?�@��          >  >  ?� �  �������� ~       � �          0���/�  `  ?��     ? �  ���� 0               ?� �  >          �       � �          >���/�  �  ��     ? ~   ���� �          ?    ?� �  � #���� �  � ?� � �          0������ `  #� ?������   ����� � 0               >> �  "            �     �          ?��������  � ?������ �  ��������          ?   ?� `  � >�� �  � ?��� �          8���?� `  "� "   ���� 0              >> �  "            �    �          ?���?���  � " �  ��|���          ? 8�?� `  � " �  �?��� �          8�����  `  #� >��    �����  0           8   >> �  "            �    �          ?ǔ����  � >�� �  ���x?���          ? |>��� `  � >�� �  �>�_� �          8�����!� `  "� "   ���a� 0           |  ?� �  "            �>  � �          ?���rB!��  � " �  ��`�9!��          ?�|��� `    �� ��   �  �>��� 0          <������ `  #   �  �   �����A 0          �|  � �  "� "   �> �� �          ?����R ��  � >�� �  ����A�          ?�|  �� `     �  � �  �> �G� 0          <���� `  "            ���`� 0          �|  � �  "� #����   �>  � �          ?����@�  � #���� �  ���a ��          ?�8   � `    �� ��   �  �   � 0          >C���� `  #   �  �   !��A� 0          �8   � �  "� "    �   � �          ?�C�����  � >�� �  �!��A��          ?�    � `     �  � �  �    � 0          > ����� `  "             A��A��0          �    � �  "� #����    �    � �          ?�������  � #���� �  �A��A���          ?�       8`             �  �       0          ?���?�  `  #   �  �   ����A�  0           �       ?�  "�           p       �          ?����?� ?�  � < �  � �  ����A� �          ?�       8�    ������ �  �       p          ??��?�  �  "  """""    ���A�  p           �       ?   "� -������    p       �          ?�?��?� ?�  � /������ �  ���A� �          ?�      ��             �  �     � xp          ?� }܂�  �  #           ��>�A�� p           x       �   "� /������    <       �          ?� }܂� ��  � ?������ �  ��>�A��          ?�       ��  ?������A�  �       pp          ?� a��� �  ";�����}�  ��0��C�� p           8       �   "� wwwwwP �          �          ?� a�����  �/������A�  ��0��C���          �  8   ��         A `  �      �`          � A���� �  #;�     '}�  �� �qO�� `           <  8   �   "��������<��         ��          � A������  �?������A�  �� �qO����          �  |   ��  ?������A�  �  >   ��          � ��?���  "+�"""""}��  �  �I�� �             |   �   "��������<�P     >   �           � �������  �/������A�  �  �I_����          �� �   �  �0     pA�  ��    ��          �  �|�@�  #��     tA�  �  �I�`  �           � �   �   "  ������  P   �    �           �� �|�O��  �?������A�  �� �I�`'��          �� �   �  ������A�  ��    ��          � �p� �  #���������}��  �  �I�`  �           � �   �   "  wwwww@  P   �    �           ���p���  �������A�  �� �I�`��          �� �   >�  ������A�  ��    �          �  `� �  #���������}��  �  � �` �           � �   ?�   "           P   �    �           �� `�?��  �������A�  �� � �`��          �� |   |�         A�  �� >   >�          �  @� �  #���     ?}��  �  � �` �           � |   �   "           P    � >   ?�           �� @���  �      8A�  �� � �`?��          �| 8  ��  �x��A�  �>    ��          � �� �  #�������}��  �  � �@ �           � 8  ��   "	� �x�<�P    �    ��           �������  �������A�  �� � �@���          �    �   ������A�  ���   ��          �   �    #����H��}��  �� � �@ �            �    ��   "	�      <�P    �   ��           ��  ���   ��H��A�  ���� �C���          ���   �    �x� A�  ���   ��          ��  ��    #�������|Ax�  ��   �@ �            �   ��   "       � P    ?�   ��           ��� ����   �������A�  ���  �G���          ���   ?     �x� A�  ���   ��          ��  �     #����x�}��  ��   �  �            �   ?��   "  ����  P    ?�   ��           ��� �?��   �������A�  ���  ����          ��  �           A�  ��?� �            ��         #���������}��  ��                   ?�  ���   "           P    �� ���           ���  ���   �   ���A�  ���� ���           ��  �p          A �  ��?� �8           ��     p   #���������}�  ��     8             �  ���   "          P    �� ���           ���  ���   �   ���A �  ���� ���           ��� ���>          A �  ��� ��           ��    �>   #���������}�  ��    �             �� ��?�   "	�      <�P     �� ��           ���� ����   �I$���hA�  ���� ���           ������<          A �   ��������           ��   �<   #���������}�   ���   �             �����   "	�      <�P    ?����?�           ���������   �   ���A �   ���������           ������< |          A �   ����� >           ���   < |   #��������A   ���    >             ������   "              ������           ���������   �   ���A �   ���������            ��  � �          A �   �?� � |            ��  � �   #���������}�   �?� � |             �����    "              �����            ���������   �I$���hA�   ��������            �� ��          A �   ?�� ?� �            �� ��   #���������}�   ?�� ?� �             ���?�    "              ����             ��������   �   ���A �   ?��������            � ��� �          A �   ?� �� �            � ��� �   #���������}�   ?� �� �             �  ��    "               �� ��             ��������   �   ���A �   ?��������            ?� �� �          A �   ���� �            ?� �� �   #���������}�   ���� �              �� ��    "	�      <�     � ?��             ?��������   �I$���hA�   ��������            ��    �          A �   ��    �            ��    �   #���������}�   ��    �              �����    "	�      <�     ?�����             ��������   �   ���A �   ��������            ��    ?�          A �   ��    �            ��    ?�   #��������A   ��    �              �����    "               �����             ��������   �   ���A �   ��������            ��    �          A �   ��    ?�            ��    �   #���������}�   ��    ?�              �����    "               �����             ��������   �I$���hA�   ��������            ��   �           A �   ��    ��            ��   �    #���������}�   ��    ��              ����     "               ����              �������    �   ���A �   ��������            ��   �           A �   ��   �             ��   �    #���������}�   ��   �               ����     "                ����              �������    �   ���A �   �������             ���  �           A �    ���  �             ���  �    #���������}�    ���  �                ?���     "	�      <�      ���              �������    �I$���hA�    �������              ��  ��           A �    ?��  �              ��  ��    #���������}�    ?��  �                ��      "	�      <�      ���               ������    �   ���A �    ?������              ?�����           A �    �����              ?�����    #��������A    �����                 �      "                 ?�                ?������    �   ���A �    ������              ������           A �    ������              ������    #���������}�    ������                         "                                   ������    �I$���hA�    ������              �����            A �    ������              �����     #���������}�    ������                         "                                   �����     �   ���A �    ������              �����            A �    �����               �����     #���������}�    �����                          "                                   �����     �   ���A �    �����                �����            A �     ����                �����     #���������}�     ����                          "	�      <�                          �����     Bm��rI$�A
�     ����                ?����            A �     ����                ?����     #���������}�     ����                          "	�      <�                          ?����     ���   A�     ����                ���             A �     ����                ���      #��������A     ����                          "                                    ���      ���   A�     ����                 ���             A �      ��                  ���      #���������}�      ��                           "                                     ���      Bm��rI$�A
�      ��                  ��             A �      ��                  ��      #���������}�      ��                           "                                     ��      ���   A�      ��                                  A �                                    #���������}�                                    "                                              ���   A�                                           A �                    ��������������������������}�������������������  �����������������	�      <�������������������                  Bm��rI$�A
�                    ���������������       A ������������������   �              ����������}�                 �  �              �	�      <�                 �  ������������������   A������������������   ���������������       A ������������������   �              ���������A                 �  �              �                           �  ������������������   A������������������   ���������������       A ������������������   �              ����������}�                 �  �              �                           �  ���������������Bm��rI$�A
������������������   p                      A �                   ��������������������������}�������������������  �����������������          ������������������  p               ���   A�                   p                      A �                   ��������������������������}�������������������  �����������������          ������������������  p               ���   A�                   p                      A �                   ��������������������������}�������������������  �����������������	�      <�������������������  p               Bm��rI$�A
�                   p                      A �                   ��������������������������}�������������������  �����������������	�      <�������������������  p               ���   A�                   p                      A �                   �������������������������A������������������  �����������������          ������������������  p               ���   A�                   p                      A �                   ��������������������������}�������������������  �               "                          �  t���m�$�Im�ےI$�Bm��rI$�A
�I$���m�$�Im�ےI'   p                      A �                   ��������������������������}�������������������  �               "                          �  p����   ?���   ���   A�  ����   ?���     p                      A �                   ��������������������������}�������������������  �               "                          �  p����   ?���   ���   A�  ����   ?���     p                      A �                   ��������������������������}�������������������  �               "	�      <�                �  t���m�$�Im�ےI$�Bm��rI$�A
�I$���m�$�Im�ےI'   p                      A �                   ��������������������������}�������������������  �               "	�      <�                �  p����   ?���   ���   A�  ����   ?���     p                      A �                   �������������������������A������������������  �               "                          �  p����   ?���   ���   A�  ����   ?���     p                      A �                   ��������������������������}�������������������  �               "                          �  t���m�$�Im�ےI$�Bm��rI$�A
�I$���m�$�Im�ےI'   p                      A �                   ��������������������������}�������������������  �               "                          �  p����   ?���   ���   A�  ����   ?���     p                      A �                   ��������������������������}�������������������  �               "                          �  p����   ?���   ���   A�  ����   ?���     p                      A �                   ��������������������������}�������������������  �               "	�      <�                �  t���m�$�Im�ےI$�Bm��rI$�A
�I$���m�$�Im�ےI'   p                      A �                   ��������������������������}�������������������  �               "	�      <�                �  p����   ?���   ���   A�  ����   ?���     p                      A �                   �������������������������A������������������  �               "                          �  p����   ?���   ���   A�  ����   ?���     p                      A �                   ��������������������������}�������������������  �               "                          �  t���m�$�Im�ےI$�Bm��rI$�A
�I$���m�$�Im�ےI'   p                      A �                   ��������������������������}�������������������  �               "                          �  p����   ?���   ���   A�  ����   ?���     p                      A �                   ��������������������������}�������������������  �               "    x�                   �  p����   ?���   ��    A�  ����   ?���     p                      A �                   ���������������������}����}�������������������  �               "	� }�߀<�                �  t���m�$�Im�ےI$��H   [hA�I$���m�$�Im�ےI'   p                      A �                   ���������������������}����}�������������������  �               "	� }���<�                �  p����   ?���   �     ?�A �  ����   ?���     p                      A �                   ��������������������}����A������������������  �               "   }���                  �  p����   ?���   �     �A �  ����   ?���     p                      A �                   ���������������������}����}�������������������  �               "   }���                  �  t���m�$�Im�ےI$��@   hA�I$���m�$�Im�ےI'   p                      A �                   ���������������������}����}�������������������  �               "   }���                  �  p����   ?���   �     �A �  ����   ?���     p                      A �                   ���������������������}����}�������������������  �               "   +}���                  �  p����   ?���   �     �A �  ����   ?���     p                      A �                   ���������������������}����}�������������������  �               "	� +}���<�                �  t���m�$�Im�ےI$��    hA�I$���m�$�Im�ےI'   p                      A �                   ���������������������}����}����������������������               "	� +}���<�                ���p����   ?���   �     �A �  ����   ?���     p                      A �                ����������������������}����A������������������ �               "   +}���                  � p����   ?���   �     �A �  ����   ?���  ��p                      A �                �����������������������}����}������������������� �               "   +}���                  � t���m�$�Im�ےI$��    hA�I$���m�$�Im�ےI'��p                      A �             ��������������������������}����}��������������  �� �               "   +}���               ���� p����   ?���   �     �A �  ����   ?�������p                 ?��  A �             �  ���������������������������}��������������� �� �               "   +@W�               ��� p����   ?���   �  ?���A �  ����   ?�������p                �   A �             �  ���������������������������}��������������� �� �               "	� *���<�             ��� t���m�$�Im�ےI$��� �hA�I$���m�$�Im����'��p                   � A �             �  �����������������������}����}��������������� �� �               "	� (}��8<�             ��� p����   ?���   �    ��A �  ����   ?�������p                    A �             �  ����������������������}�ߟ�A�������������� �� �               "   !}�ߨ               ��� p����   ?���   �    7�A �  ����   ?�������p                     A �             �  �����������������������}����}��������������� �� �               "   #}���               ��� snI$�F�m��I$m��]�   hA��nI$�F�m��I������p                     A �             �  �����������������������}����}��������������� �� �               "   }���               ��� w�   ����   �����     �A ����   ����  ������p                @     A �             �  �����������������������}����}��������������� �� �               "   }���               ��� w�   ����   ����� @   �A ����   ����  ������p                      A �             �  �����������������������}����}��������������� �� �               "	� +}���<�             ��� snI$�F�m��I$m��]�    hA��nI$�F�m��I������p                      A �             �  �����������������������}����}��������������� �� �               "	� +}���<�             ��� w�   ����   �����     �A ����   ����  ������p                      A �             �  ����������������������}����A�������������� �� �               "   +}���               ��� w�   ����   �����     �A ����   ����  ������p                      A �             �  �����������������������}����}��������������� �� �               "   +}���               ��� snI$�F�m��I$m��]�    hA��nI$�F�m��I������p                      A �             �  �����������������������}����}��������������� �� �               "   +}���               ��� w�   ����   �����     �A ����   ����  ������p                      A �             �� �����������������������}����}������������������ �             ��   +}���  �            ~�� w�   ����   �� �     �A � ��   ����  ������p            ��       A �            � �����������������I#����}����}�I��������������� �           �I"	� +}���<�I��          y��� snI?�F�m��I$h�݂    hA� nI$�F�m��I������p  ,�        m��       A ��           � ������?����������I#����}����}�I$�������������� �  �        �I"	� +}���<�I$�          w��� w� �����   �m���     �A ��|   ����  ������p  w�        o��       A ���           � ����� ����������� #���}����A$�������������� �  ��        � "   +}���  $�          o��� w� ������   �o���     �A ���|   ����  ������p  �`        ���       A ��           � �����_���������I#����}����}�H �������������� �  ��        I"   +}���  H �          o��� snI��F�m��I$k��݂    hA��nI$�F�m��I������p  �P        m��       A ��           ������� /����������I#����}����}�I$���������������� � ��        �I"   +}���  I$�          _`� w�������   �m���     �A ��|   ����  ������p �0        m��       A ��           ��������_/����������I#����}����}�I$���������������� � ��        �I"   +}���  I$�          ^`� w�������   �m���     �A ��|   ����  ������p ��        m��       A ��           ������������������I#����}����}�I$��������������� � �0        �I"	� +}���<�I$�          ^`� snI��F�m��I$km��Bm�   �A
��nI$�F�m��I�����p �P        m��       A ��           �0�����������������I#����}����}�I$���������������� � �0        �I"	� +}���<�I$�          ~�`� w��p����   �m���     A��|   ����  ������p �p        o��       A ��           ������������������ #���}����AI$���������������� � �p        � "   +}���  I$�          `� w��p����   �o���     A��|   ����  ������p  @�        ���       A ���           � ����������������I#����}����}�$�������������� �  �`        I"   +}���  $�          ��� snI��F�m��I$k���Bm�   �A
���nI$�F�m��I������p  1�        m��       A ��           � �����_����������I#����}����}�H �������������� �  ��        �I"   +}���  H �          ��� w� ������   �m���     A��|   ����  ������p  �        l        A ��           � ������?����������������}����}�I$�������������� �  �        ���   +}���  I$�          ��� w� �����   �l �     A��|   ����  ������p                ?��  A � �           � ����������������� #��������}��$������������ �� �           � "	� +@W�<��$�          ��� snI?�F�m��I$h  Bm�?�� �A
� �nI$�F�m��I������p                �   A �             �� ���������������������������}�������������� �� �               "	� *���<���          ��� w�   ����   ������ � A�  |   ����  ������p                   � A �             �  ����������������������}����A�������������� �� �               "   (}��8               ��� w�   ����   �����   � A����   ����  ������p                    A �             �  �����������������������}����}��������������� �� �               "   !}���               ��� snI$�F�m��I$m��\Bm�   4�A
��nI$�F�m��I������p                     A �             �  �����������������������}����}��������������� �� �               "   #}���               ��� w�   ����   �����    A����   ����  ������p                     A �             �  �����������������������}����}��������������� �� �               "   }���               ��� w�   ����   �����    A����   ����  ������p                @     A �             �  �����������������������}����}��������������� �� �               "	� }���<�             ��� snI$�F�m��I$m��\Bm�   �A
��nI$�F�m��I������p                      A �             �  �����������������������}����}��������������� �� �               "	� +}���<�             ��� w�   ����   �����     A����   ����  ������p                      A �             �  ����������������������}����A�������������� �� �               "   +}���               ��� w�   ����   �����     A����   ����  ������p                      A �             �  �����������������������}����}��������������� �� �               "   +}���               ��� t���m�$�Im�ےI$�Bm�   �A
�I$���m�$�Im����'��p                      A �             �  �����������������������}����}��������������� �� �               "   +}���               ��� p����   ?���   �     A�  ����   ?�������p                      A �             �  �����������������������}����}��������������� �� �               "   +}���               ��� p����   ?���   �     A�  ����   ?�������p                      A �             �  �����������������������}����}��������������� �� �               "	� +}���<�             ��� t���m�$�Im�ےI$�Bm�   �A
�I$���m�$�Im����'��p                      A �             �  �����������������������}����}��������������� �� �               "	� +}���<�             ��� p����   ?���   �     A�  ����   ?�������p                      A �             �������������������������}����A������������������ �               "   +}���                  � p����   ?���   �     A�  ����   ?�������p                 q�  A �             ��������������������������0���}������������������� �               "   +0��                  � t���m�$�Im�ےI$�Bm�q��A
�I$���m�$�Im����'��p                m�[  A �             ��������������������������@���}������������������� �               "   (@��                  � p����   ?���   �m�[  A�  ����   ?�������p                ���� A �                �����������������������  �}������������������� �               "                        � p����   ?���   ����� A�  ����   ?���  ��p                ?}��x A �                ������������������������ ��}������������������� �               "	�  � �<�                � t���m�$�Im�ےI$�Bm�}��|�A
�I$���m�$�Im�ےI'��p                m6iP A �                ����������������������� �'�}������������������� �               "	�   � <�                � p����   ?���   �m6iP A�  ����   ?���  ��p                      A �                ���������������������������A������������������ �               "                          � p����   ?���   ���   A�  ����   ?���  ��p                      A �                ����������������������������}������������������� �               "                          � t���m�$�Im�ےI$�Bm��rI$�A
�I$���m�$�Im�ےI'��p                      A �                ����������������������������}������������������� �               "                          � p����   ?���   ���   A�  ����   ?���  ��p                      A �                ����������������������������}������������������� �               "                          � p����   ?���   ���   A�  ����   ?���  ��p                      A �                ����������������������������}������������������� �               "	�      <�                � t���m�$�Im�ےI$��I$���hA�I$���m�$�Im�ےI'��p                      A �                ����������������������������}������������������� �               "	�      <�                � p����   ?���   �   ���A �  ����   ?���  ��p                      A �                ���������������������������A������������������ �               "                          � p����   ?���   �   ���A �  ����   ?���  ��p                      A �                ����������������������������}������������������� �               "                          � t���m�$�Im�ےI$��I$���hA�I$���m�$�Im�ےI'��p                      A �                ����������������������������}������������������� �               "                          � p����   ?���   �   ���A �  ����   ?���  ��p                      A �                ����������������������������}������������������� �               "                          � p����   ?���   �   ���A �  ����   ?���  ��p                      A �                ����������������������������}������������������� �               "	�      <�                � t���m�$�Im�ےI$��I$���hA�I$���m�$�Im�ےI'��p                      A �                   ��������������������������}����������������������               "	�      <�                ���p����   ?���   �   ���A �  ����   ?���     p                      A �                   �������������������������A���������������������               "                          ���p����   ?���   �   ���A �  ����   ?���     p                      A �                   ��������������������������}����������������������               "                          ���t���m�$�Im�ےI$��I$���hA�I$���m�$�Im�ےI'   p                      A �                   ��������������������������}����������������������               "                          ���p����   ?���   �   ���A �  ����   ?���     p                      A �                   ��������������������������}�������������������  �               "                          �  p����   ?���   �   ���A �  ����   ?���     p                      A �                   ��������������������������}�������������������  �               "	�      <�                �  t���m�$�Im�ےI$��I$���hA�I$���m�$�Im�ےI'   p                      A �                   ��������������������������}�������������������  �               "	�      <�                �  p����   ?���   �   ���A �  ����   ?���     p                      A �                   �������������������������A������������������  �               "                          �  p����   ?���   �   ���A �  ����   ?���     p                      A �                   ��������������������������}�������������������  �               "                          �  snI$�F�m��I$m��]�I$���hA��nI$�F�m��I$m��   p                      A �                   ��������������������������}�������������������  �               "                          �  w�   ����   �����   ���A ����   ����   ���   p                      A �                   ��������������������������}�������������������  �               "                          �  w�   ����   �����   ���A ����   ����   ���   p                      A �                   ��������������������������}�������������������  �               "	�      <�                �  snI$�F�m��I$m��]�I$���hA��nI$�F�m��I$m��   p                      A �                   ��������������������������}�������������������  �               "	�      <�                �  w�   ����   �����   ���A ����   ����   ���   p                      A �                   �������������������������A������������������  �����������������          ������������������  p               �   ���A �                   ���������������       A ������������������   �              ����������}�                 �  �              �                           �  ����������������I$���hA������������������   ���������������       A ������������������   �              ����������}�                 �  �              �                           �  ����������������   ���A ������������������   ���������������       A ������������������   �              ����������}�                 �  �              �                           �  ����������������   ���A ������������������                          A �                    ��������������������������}�������������������  �����������������	�      <�������������������                  �I$���hA�                                          A �                   ��������������������������}�������������������  �����������������	�      <�������������������                  �   ���A �                                          A �        �          �������������������������A�����������������  �����������������          ������������������                  �   ���A �                             ?�            A �        �          �������������������������}����������?��������  �����������������          ������������������          @      �I$���hA�                           ?�            A �        �          �������������������������}����������?��������  �����������������          ������������������          @      �   ���A �                      �  ?�            A �    �  �          ������������������������}���������?��������  �����������������          ����������������         a`     �   ���A �      �0�0               �  ?�            A �    �  �          ������������������������}���������?��������  ����������������	�      <�������?����������        �a `     Bm��rI$�A
�      �0�0               �  �            A �    �  �          ������������������������}���������?��������  ���������������	�      <�������?����������        �� `     ���   A�      �p�0               �              A �    �            ������������������������A�����������������  �������?\�������          �������w���������        ���     ���   A�      �Q�p               �               A �    ��            �������������������������}������������������  �������?�������          ����������������       A�� �     Bm��rI$�A
�     ��qp               �   �           A �    �   |         ������������������������}������������������  ������>=�������          ������ߏ�������       #���@�     ���   A�    ��a p�              ?�=x�           A �    �� �               ��    #���������}�      ��@s@              ><=x�    "              � �              �����    ���   A�     ����s@              �}p�           A �    �>��               ႏ�    #���������}�      ��G�              �}p�    "	�      <�    �>��               ����    Bm��rI$�A
�     ����              ���           A �    �X��             �O�`    #���������}�    ����0              � ��    "	�      <�    � X��             ����`    ���   A�    ����0              �  �           A �    � ���             8�O��    #��������A    �ç�H              �   �    "              �   �             8�O��    ���   A�    ��'�X              �  �           A �    �  ��             |�G�H    #���������}�    >��#�$              �   �    "              �   �             |�G�x    Bm��rI$�A
�    >��#�<                 �           A �     �  ��            ~��G� �   #���������}�   ?a��#� |                �    "               �  �            ��G�0�   ���   A�   ?���#�|              >  w�           A �     �  ;��            ~������   #���������}�   �p��a�D              >  �    "               �  ��            ���È�   ���   A�   ����a�D               >  ��           A �        }�             ~qɜ��     #���������}�    �8��C�                 6  �    "	�      <�        �             ~q���     Bm��rI$�A
�    �8��C�                 >  ��           A �        |�             �����     #���������}�   ?����G�                 >  �    "	�      <�        �             ����     ���   A�   ?����G�                   ��           A �        |             ���     #��������A   ?���č�                   8�    "                               �㉛8    ���   A�   ?����͜               �  p           A �     p  8�            �����    #���������}�    �������                      "                  �            ��ӑ�    Bm��rI$�A
�    ������߀             �              A �   � �   �             ����p    #���������}�    ~�����                       "             �     �             ���    ���   A�    ~�����             �   �          A �   ��   �             �����    #���������}�    ~��цp               @   �   "             �     �            �G����   ���   A�   ~#�цq�            ?�   q�          A �   ��   8�             ��� ��    #���     ?}�    ?����~�             ?  �   q�   "	�������<�   � P   8�             q��� ���   Bo������A
�   8�S��~��            >�   ��   ������A �   ��   |p             ���'�     #���"""""=}�    ?�����             >  @   ��   "	�������<�         |p            0`�G�'� �   ������A�   0~#���p            x�  �           A �   <��   �              ����S�   #��     <A    ?��܏�)�            x    �    "  ������    <     �             xd���S�   ������A�   <2���)�              �  �                     �p   �            �w���   �������������   ;����                   �   �������������          �            �h�� 8  �������������   4?���            �    �8  �������������   p     �            �=���S    A � �   �����)�            �     �8  ��߾���~���}�   p      �            ��?���S8  �������������   q�����)�           �   � �  �������������   �   � |            ������   A � �   ������           �      �  ��߾���~���}�   �      |           �����|�  �������������   ����>��           �   � p                   �   � 8            �������  �������������    ������           �      p  �������������   �      8           �����<��  �������������   ������           �  ��    �������������  �  ��              ;����w��    A � �@   ���;��           �  �     ߾���~���}��  �  ��             ����9w��  �������������  �������           �  ��   �������������  �  ��  �            ?�����     A � �@   ����            �  �    ߾���~���}��  �  �   �           ���� 0�  �������������  ��� �             8� �                  � �� À           �����   �������������   �k����             (�  �  �������������  � �  À          ��� `�  �������������  ��c�0���            |�   �������������  � >�  ��           ��ҟ���    A � �   �~�O���               �    ��߾���~���}�  �  �   ��          �ҟ���  �������������  ��@�O����            �� >   �������������  � �  �            �}�����   A � �    ~>�����             ��     ��߾���~���}�  � A�   �           ������  �������������  �~ �����           ��  �                 � � ?��            �������  �������������    |�����            �  � �������������  � �  �           �����ǀ �������������  �|�����             ��  � �������������     � ?��          �������    A � �@  ��w��?��              (�  � ߾���~���}��     �  �          ��9���� �������������  ������            �    � �������������       ?��          0�}ܿ���    A � �@  �>�_�?��             �    � ߾���~���}��    I    �          >�ܿ���� �������������  ��_���            |   > �                   >     �           ��������  �������������  ������                   � �������������           �          .��������� �������������  �A������            8   � �������������      �  �          @l������   A � �   �K����             (     � ��߾���~���}�          �          N|������� �������������  '�C����              �� � �������������      ��  �          |�ȟ��@  A � �  >O�O��                #� � ��߾���~���}�       �  �          |�Ȝ\�� �������������  >O�N.��             w� �                  �   �� �           ��G���@ �������������   ?��#��               w� � �������������   �   ;� �           ��F���� �������������   ?��#D��          �   /� �   A � �@  �   � �           ��y��p@   A � �@   ?��<�p8           �   /� � ߾���~���}��  �   � �           ��y��s� �������������   ?��<�p9�             � �   A � �@   �  � �          ����� @   A � �@  ��?�@�               � � ߾���~���}��   �   � �          ������ �������������  ��?�@��          >  >  ?� � �������������      � �          0���/�  `                 ���� 0               ?� � �������������       � �          >���/�  � �������������  ���� �          ?    ?� �  A � �  � ?� � �          0������ `  A � �  ����� � 0               >> � ��߾���~���}�  �     �          ?�������� �������������  ��������          ?   ?� `  A � �  � ?��� �          8���?� `  A � �  ���� 0              >> � ��߾���~���}�  �    �          ?���?��� �������������  ��|���          ? 8�?� ` �������������  �?��� �          8�����  `                  �����  0           8   >> � �������������  �    �          ?ǔ���� �������������  ���x?���          ? |>��� `   A � �@  �>�_� �          8�����!� `   A � �@  ���a� 0           |  ?� � ߾���~���}��  �>  � �          ?���rB!�� �������������  ��`�9!��          ?�|��� `   A � �@  �>��� 0          <������ `   A � �@  �����A 0          �|  � � ߾���~���}��  �> �� �          ?����R �� �������������  ����A�          ?�|  �� ` �������������  �> �G� 0          <���� `                 ���`� 0          �|  � � �������������  �>  � �          ?����@� �������������  ���a ��          ?�8   � `  A � �  �   � 0          >C���� `  A � �  !��A� 0          �8   � � ��߾���~���}�   �   � �          ?�C����� �������������  �!��A��          ?�    � `  A � �  �    � 0          > ����� `  A � �   A��A��0          �    � � ��߾���~���}�   �    � �          ?������� �������������  �A��A���          ?�       8` �������������  �       0          ?���?�  `                 ����A�  0           �       ?� �������������   p       �          ?����?� ?� �������������  ����A� �          ?�       8�   A � �@  �       p          ??��?�  �   A � �@  ���A�  p           �       ?  ߾���~���}��   p       �          ?�?��?� ?� �������������  ���A� �          ?�      ��   A � �@  �     � xp          ?� }܂�  �   A � �@  ��>�A�� p           x       �  ߾���~���}��   <       �          ?� }܂� �� �������������  ��>�A��          ?�       �� �������������  �       pp          ?� a��� �                 ��0��C�� p           8       �  �������������          �          ?� a����� �������������  ��0��C���          �  8   ��  A � �  �      �`          � A���� �  A � �  �� �qO�� `           <  8   �  ��߾���~���}�         ��          � A������ �������������  �� �qO����          �  |   ��  A � �  �  >   ��          � ��?���  A � �  �  �I�� �             |   �  ��߾���~���}�     >   �           � ������� �������������  �  �I_����          �� �   � �������������  ��    ��          �  �|�@�                 �  �I�`  �           � �   �  �������������   �    �           �� �|�O�� �������������  �� �I�`'��          �� �   �   A � �@  ��    ��          � �p� �   A � �@  �  �I�`  �           � �   �  ߾���~���}��   �    �           ���p��� �������������  �� �I�`��          �� �   >�   A � �@  ��    �          �  `� �   A � �@  �  � �` �           � �   ?�  ߾���~���}��   �    �           �� `�?�� �������������  �� � �`��          �� |   |� �������������  �� >   >�          �  @� �                 �  � �` �           � |   �  �������������    � >   ?�           �� @��� �������������  �� � �`?��          �| 8  ��  A � �  �>    ��          � �� �  A � �  �  � �@ �           � 8  ��  ��߾���~���}�    �    ��           ������� �������������  �� � �@���          �    �   A � �  ���   ��          �   �    A � �  �� � �@ �            �    ��  ��߾���~���}�    �   ��           ��  ���  �������������  ���� �C���          ���   �  �������������  ���   ��          ��  ��                   ��   �@ �            �   ��  �������������    ?�   ��           ��� ����  �������������  ���  �G���          ���   ?                   ���   ��          ��  �     <          �  ��   �  �            �   ?��   <          �    ?�   ��           ��� �?��                  ���  ����          ��  �                   ��?� �            ��         <          �  ��                   ?�  ���   <          �    �� ���           ���  ���                  ���� ���           ��  �p                  ��?� �8           ��     p   <          �  ��     8             �  ���   <          �    �� ���           ���  ���                  ���� ���           ��� ���>                  ��� ��           ��    �>   ?������������  ��    �             �� ��?�   >          �     �� ��           ���� ����   �����������   ���� ���           ������<   �����������    ��������           ��   �<   >          �   ���   �             �����   >          �    ?����?�           ���������                   ���������           ������< |     ����   �   ����� >           ���   < |   #�����������   ���    >             ������   "              ������           ���������   ������������   ���������            ��  � �   ��������   �?� � |            ��  � �   "       �?� � |             �����    "              �����            ���������        �   ��������            �� ��        �   ?�� ?� �            �� ��   #�������   ?�� ?� �             ���?�    "              ����             ��������   ��������   ?��������            � ��� �   ��������   ?� �� �            � ��� �   "       ?� �� �             �  ��    "               �� ��             ��������        �   ?��������            ?� �� �     �� ��   �   ���� �            ?� �� �   #��� �  ���   ���� �              �� ��    "         � ?��             ?��������   ��������   ��������            ��    �   ��� �  ����   ��    �            ��    �   "             ��    �              �����    "  ����       ?�����             ��������     ����   �   ��������            ��    ?�     �� ��   �   ��    �            ��    ?�   #��� �  ���   ��    �              �����    "         �����             ��������   ��������   ��������            ��    �   ��� �  ����   ��    ?�            ��    �   "             ��    ?�              �����    "  ����       �����             ��������     ����   �   ��������            ��   �               �   ��    ��            ��   �    #��� �  ���   ��    ��              ����     "               ����              �������    ��� �  ����   ��������            ��   �    ������������   ��   �             ��   �    "             ��   �               ����     "                ����              �������               �   �������             ���  �               �    ���  �             ���  �    #�����������    ���  �                ?���     "                ���              �������    ������������    �������              ��  ��    ������������    ?��  �              ��  ��                    ?��  �                ��                        ���               ������    ������������    ?������              ?�����    ������������    �����              ?�����                    �����                 �                         ?�                ?������    ������������    ������              ������    ������������    ������              ������                    ������                                                              ������    ������������    ������              �����                      ������              �����     ?������������    ������                         ?������������                         �����                      ������              �����                      �����               �����     ?������������    �����                          ?������������                         �����                      �����                �����                       ����                �����     ?������������     ����                          ?������������                          �����                       ����                ?����                       ����                ?����     ?������������     ����                          ?������������                          ?����                       ����                ���                        ����                ���      ?������������     ����                          ?������������                          ���                        ����                 ���                         ��                  ���      ?������������      ��                           ?������������                           ���                         ��                  ��                         ��                  ��      ?������������      ��                           ?������������                           ��                         ��                                                                            ?������������                                    ?������������                                                                                                                                      ?������������                                    ?������������                                                                                                                                      ?������������                                    ?������������                                                                                                                                      ?������������                                    ?������������                                                                                                                                      ?������������                                    ?������������                                                                                                                                      ?������������                                    ?������������                                                                                                                                      ?������������                                    ?������������                                                                                                                                      ?������������                                    ?������������                                                                                                                                      ?������������                                    ?������������                                                                                                                                      ?������������                                    ?������������                                                                                                                                                                         