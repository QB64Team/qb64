��b  �-               �     �                            �     �                            �     �                            �     �                           �     �                           �     �                           �     �                           �     �                           �     �                           �     �                           �     �                           �     �                          ��y���6�<�                          ��y���6�<�                          ��y���6�<�                          ��y���6�<�                          �l��6ݳf�                          �l��6ݳf�                          �l��6ݳf�                          �l��6ݳf�              ����������� ��}�͘?ٿ~�  ���������������������� ��}�͘?ٿ~�  �����������            ��}�͘?ٿ~�                          ��}�͘?ٿ~�                                                                                                      ��Ͷ͘?ٰ`�                                                                                                                                            �lͶ͘��f�                                                                                                                                            ��}�����<�m�                                                                                                                                                                                                                                                                                                      �                                                         