��]  Ta�                                                                         ������������������������������������                                                                                                            ������������������������������������                                    ������������������������������������                                    ������������������������������������                                    ������������������������������������                                    ������������������������������������                                     ?����������                        ��         ?������������������������ ?����������                                                            ������������������������������������                                    ������������������������������������                                     ?����������                   ���� ��0       ?�������������������   � ?����������                   ����   0                                ������������������������������������  0 0  �                         0  ������������������������������������  0 0  �                             ?����������                   ���� ��0 0  �   ?�������������������  8� ?����������                   ����   0 0  �                            ������������������������������������  7�;�<���                    ��  �������������������������������� ��  7�;�<���                          ?����������                   ���� ��7m�3f͛��?���������������������� ?����������                   � �   7m�3f͛��                         ��ə�̟2d���������������������������                               ��  ��������������������������������  ��                                     ?ɜ�̟2d��                   ���� ��         ?���������������������� ?����������                   � �                                     ��ɒLș2d�?�������������������������                               ��  �������������������������������� ��                                     ?ɘ��Ó��                   ���� ��         ?�������������������  8� ?����������                   ����                                     ������������������������������������                                 0  ������������������������������������                                     ?����������                   ���� ��         ?�������������������   � ?����������                   ����                                     ������������������������������������                                    ������������������������������������                                     ?����������                        ��         ?������������������������ ?����������                                                            ������������������������������������                                    ������������������������������������                                    ������������������������������������                                    ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������?����������?������������                                                                                                            ���������������﮿�����������������                                                                                                            ���������������ﯿ����������������                                                                                                            ����Î?�m��go�������g��e����                                                                                                            ���w�u���6��q�[����6����k�u����                                                                                                            ���w�����������[����������-����                                                                                                            ���w�}�����������[�/�������?�����                                                                                                            ���w�u�������[�.�������k�u����                                                                                                            ����Î��n��u��]�����u�ߜm����                                                                                                            ������������������������������������                                                                                                            ������?�����������������������������                                                                                                            ������������������������������������                                                                                                            �����������������������������������                                                                                                            ����������������������������������                                                                                                            ����������������������������������                                                                                                            ���?q��?���f3���q�?�8~8�s����U���                                                                                                            ���~鮮��u�k����������]u�u���U���                                                                                                            ���~����u�k����������~��u���U���                                                                                                            ���~�����u�k���������u�}��{u���U���                                                                                                            ���~뮮��u�k���n�����u�}�]u�u�������                                                                                                            ������?��lv7��p�?��~�s��������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ����������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ���8�>��8���3�2Ɵ�|��3i��lq�����                                                                                                            ���u�}~���}u���uֺo��������������                                                                                                            ���u�a~���}uT��������.��(/�����                                                                                                            ���u��~����uU��}������������������                                                                                                            ���u�]~���}v���uֺ�������뫮�����                                                                                                            ���8�~������7�:������7n�lq�����                                                                                                            ���}��������������������������������                                                                                                            ���}��������������������������������                                                                                                            ������������������������������������                                                                                                            �����������������������������������                                                                                                            �������������������o���������������                                                                                                            �������������������o���������������                                                                                                            ��Ì��v�kjp�i�N1?��)�qƟ�68��q���                                                                                                            ��������������5����f���o���Z�ٮ���                                                                                                            ��݅����������t��]n�0�����۠���                                                                                                            ���u����������u���]n��������ۯ���                                                                                                            ���u������k����u����n������Z�ۮ���                                                                                                            ��Å��{�k���n�v6�����p���68������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������W�����������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ��Ì�mWÏ�����q��v���Ƨ�9�&?��                                                                                                            �����mW�w�u�]����[�����ֺ�����                                                                                                            ��݅�UW��u�]����[�����{������                                                                                                            ���u�UW��u�����[���﻽�������                                                                                                            ���u��W�w�u�]���[����ֺ�����                                                                                                            ��Å߻WÏ�������{���ƻ�9��?��                                                                                                            ������������������������������������                                                                                                            �����������������������������������                                                                                                            ������������������������������������                                                                                                            ����������o������������������������                                                                                                            ����������_�������������������������                                                                                                            ����������_�������������������������                                                                                                            ���������O�|��3i�����������������                                                                                                            ���}��]�}_�����������������������                                                                                                            ���}��]�a_�����.�����������������                                                                                                            ���}���]�]_�������������������������                                                                                                            ���}��]�]_�����������������������                                                                                                            ���~����a_����7n�����������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            �����������������������������������                                                                                                            �����������������������������������                                                                                                            �����������������������������������                                                                                                            ����8��~�~��L63?ln�j�
�i�N?���                                                                                                            �����M�k�껾��u����k��j�����5����                                                                                                            ���]�]��>�x>��u���k�����>�X.�t���                                                                                                            ���]���������u�����k�������[��u����                                                                                                            �����]���۾��u���뿛��ھ�뻮�u����                                                                                                            ��������~�~�㍴6;?�r�ھ�n�v?���                                                                                                            ������������������������������������                                                                                                            ����������������������������������                                                                                                            ������������������������������������                                                                                                            ���������������������}������������                                                                                                            ���������������������}������������                                                                                                            ���������������������}������������                                                                                                            ���N4��q�~��q���8~8a�Q?���������                                                                                                            ���7�]w۾龚뾶�������]���k��������                                                                                                            ���v_۾����>����~]��߻��������                                                                                                            ���u�_۾�������u�}�]���ۯ�������                                                                                                            ���u�]w۾뮺뾶����u�}�]���k.������                                                                                                            ���vc����~��q����~a��ߜ��������                                                                                                            ������������������������������������                                                                                                            �����������������������������������                                                                                                            ������������������������������������                                                                                                            ��������������������� �������������                                                                                                            ������������������u���������������                                                                                                            ������������������u���������������                                                                                                            ����p�js%N���3����J'�Ɵƛo����                                                                                                            ����k�����mu5�u�]m���������o�ko����                                                                                                            ���h?����muu��_w�����������o����                                                                                                            ����k�����muu�}��{����������o����                                                                                                            ����k�����muu�u�]m��������������                                                                                                            ���l��k��v������Z����������                                                                                                            �����������������������������������                                                                                                            �������������?��������������������                                                                                                            ������������������������������������                                                                                                            �����������������������������������                                                                                                            ����������������������������������                                                                                                            ����������������������������������                                                                                                            ��Ï��������~4�bq�g�c��2g����                                                                                                            ���w�u�]���ku����[�����}uw������                                                                                                            ����u�]��
�����[�����a|�v�����                                                                                                            ����u������}����[�����]}u������                                                                                                            ���w�u�]����u����[�����]u�u������                                                                                                            ��Ï����
���~7\m��o�a��g_����                                                                                                            ����������������������������������                                                                                                            �����������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                                                                                            ������������������������������������                                    