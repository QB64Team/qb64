��`  2a        �0                            �0                            �0                            �0                            �0         �                  �0         �                  �0         �                  �0         �                   0         �                   0         �                   0         �                   0         �                  3ǜ�<�}�3���                3ǜ�<�}�3���                3ǜ�<�}�3���                3ǜ�<�}�3���                ��l��3�͛6`�ٳ                ��l��3�͛6`�ٳ                ��l��3�͛6`�ٳ                ��l��3�͛6`�ٳ                 ߷��?>�͙���ٿ                 ߷��?>�͙���ٿ                 ߷��?>�͙���ٿ                 ߷��?>�͙���ٿ                                                                                   �6�0f�͙� �ٰ                                                                                                                   ٶl��3f�͘�`Ù�                                                                                                                   �3ǌ�>�}���cm�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     �                 �          �                 �                                                                            (�                 (�          *�                 *�          �                 �           �                  �         !���                 =��         ���                 ?��         -\�                 �          \�                 �        h �                  �        ����                ���        w�                 �          �                  �       �  8                           &���               ����       ��                              �                              ��@&S.                 &S        I��9��              ��9��       �x@&$                 &           P$                  P       !�� fs7                 fs0      i� y���            �� y��      -� &!                 &        H   p!                  p      �  ` 3�                ` 0     �x  ���           ��  ��     w�  �                  �          @                  @     �  ��=�               ��<    &�  ����          ��  ���    ��  � <�               � <     �  � <�               � <    ��@  � >�               � >    I��  ����          ��   ����   �x@  � ~                � ~        � >                � >   !��   ���`               ���   i�   � ~�         ��    � ~�  -�   ���@               ���    H    � >@               � >  �    �p?p               �p?  �x    ��P        ��     ��� w�    �w��               �w�        �                 �   �     ���               ���&�     � ?�       �      � ?� ��     ��Ϡ               ��π �     � �               � ��@     �x�       �      �x���     ���       �      ����@     ?w��       �      ?w��        �       �        ��      �8K�       �      �8K��      �X��       �      �X���      W�W�       �      W�W��       �       �       ��      !8��0       �      !8�� _      !D�4       _      !D�0�      ����       �      ����_        �         _        �  ?��     }�       ?��     }� ?��            ?��     ?��     >����       ?��     >����?��               ?��        ?��     >q�       ?��     >q� ~�     F       ~�     F?��     <����       ?��     <����>�               >�         �      ��       �      ��         ,p�               ,p���     =��]�       ��     =��]�         p                  p        
���             
�����      ��       ��      ��|�     =��}�       |�     =��}�         �                 �          ��L               ��@      ��             �����     =��}�       ���     =��}�         �                  �  ���     
���       ���     
�����`     ��       ��`     ��  �     =��}�         �     =��}�         �                  �  ���     ��       ���     �� ���     ,p�       ���     ,p�p�     =��]�       p�     =��]�  �      p          �      p  ���     :q�       ���     :q� ��`     F       ��`     F  �     =����         �     =����                               ���     �       ���     � ���            ���           >����             >����                                �      !=�        �      !=� �      !E8       �      !E0x��     ����       x��     ����                                        ��{�               ��{��      ����       �      ����|�     WW�       |�     WW�         �                �        �p�               �p�A�@     ���       A�@     ���>�     w��       >�     w��          �                 �?��     ��`       ?��     ���?��     � �       ?��     � �?��     ���        ?��     ���?��     �         ?��     � ��      �x?�       �      �x? _      ��?�       _      ��?��      �w�        �      �w� _      �         _      �  �      �8��       �      �8� �      �X�`       �      �X���      �?�       �      �? �      �>        �      �> �B     ��       �      �~ ��     ��       �      ���Z     ����       �      ��� �      � |�       �      � ~  o��   ���                ���  u�)    ����       ��     ���  �ր   ��                ��  �     ��                ��  [��    ��                 ��  �mJ@   ��         ?���    ��   C���   ���                 ���   )     ��                 ��    ���  ?��                 ?��   �[R�  ?��          ���   ?��    ��h  ?��                 ?��     J@   ?߀                 ?��     5��B ��                 ��     {�Ԥ ��            ��� ��     ;�Z �                 ��      �  �                 ��      o��3�                 �       ��)JR�              ����ݰ      �ֵ�@                 �        �   @                 �        [���                            �mj߀               ����        C��r                             )JR                              ֵ�                             �{�                  �          �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �                �                                                                                                                             �`                                                                                                                             �`                                                                                                           ���v��            ��p>��                                                                                                        �m�3f͘            ��`f͛0                                                                                                        3�3fy�            ��`f���                                                                                                        6m�3fy�            ̓`f��                                                                                                         6m�3f1�            ͛`f�c0                                                                                                        �3�f0�            ��0>�a�                                    