��X  .p@                                                                                                                                                                                                                �                                            �                                            �                                                                                         ��                                           ��                                           ��                                                                        �    �          ��                          �    �          ��                          �    �          ��                                                                       �   �         ���                         �   �         ���                         �   �         ���                                                                       �   �          ��                         �   �          ��                         �   �          ��                                                                       �   �          ��                         �   �          ��                         �   �          ��                                                                       �   �          ��                         �   �          ��                         �   �          ��                                                                       �   �         > ��                         �   �         > ��                         �   �         > ��                                                                       �   �         < ��                         �   �         < ��                         �   �         < ��                                                                        �    �         |  �                          �    �         |  �                          �    �         |  �                                                                                       |  @                                         |  @                                         |  @                                                                                       x >                                           x >                                           x >                                                                                         � >                                           � >                                           � >                                                                                         � ~                                           � ~                                           � ~                                                                                      � |                                        � |                                        � |                                                                           >           �?��                            >           �?��                            >           �?��                                                                   ?  `  `      �����                     ?  `  `      �����                     ?  `  `      �����                                                                  �� | x�� x      �����                    �� | x�� x      �����                    �� | x�� x      �����                                                                  �� � ��� �      ������                    �� � ��� �      ������                    �� � ��� �      ������                                                                  ��� ��� �     �������                     ��� ��� �     �������                     ��� ��� �     �������                                                                   ��� �� ��  ������                     ��� �� �  ������                     ��� �� � �  ������                                 �                                ���?��  ���x��                     ���?���  ���x��                     ���?���  ���x��                                 �                                ?���|�#� �πx �                     ?���|��  �πx �                     ?���|��� �πx �                                 ��                               >|��>���*� �� x �                     >|��>����  �� x �                     >|��>����� �� x �                                 ��                                           %�`                                           ��                               >�����=���?�� ?�� x �                                 ?��                                           d�p                                           ��                               }���������� � x                                   ��                                           ��@                                           ���                               ���������� �| x>                                   ���                                           ��8                                           ��                               ��������������x x<                                   ���                                          ��8                                          ��                               ��������������>� �< >                                 ���                                           ��                                          ���                              ���� �����>� �| <                                 ���                                           ��(                                          ���                              ��������� �x |                                 ���                                          ��(                                           ��                              ���������}��� |                                 ���                              ���>��>o�(����� �                                  ���                              ���>��>�������� �                                 ���                              �� <��<��0 ���� �                                  O��                              �� <��<��� ���� �                                 ���                              �� |� |��h?�����                                 o��                              �� |� | ���?�����                                 ���                              ��> x� x�P>�����                                 ?��                              ��> x� x ���>�����                                 ���                              ��> �� � aB�|������  @@<��  8  @             ��          �  @@<��  8  @��> �� � ���|�����                                  ���         �  @@<��  8  @�?�| ��> � ��|�����    ABAQ  D                ��0             ABAQ  D   �?�| ��> � ��|�����                                  ���             ABAQ  D   �? | ��> � �x���    A@@Q  @                M�              A@@Q  @   �? | ��> � ��x���                                  ��             A@@Q  @   ?  ���<� =� ��?��<KOY�@@Q($9�@��V                       <KOY�@@Q($9�@��V?  ���<� ?����?��                                  ?��         <KOY�@@Q($9�@��V> ~ �� |� ��ǀ~���JQe@@$Q($E9QY              �         �JQe@@$Q($E9QY> ~ �� |� � �ǀ~��                                  ��         �JQe@@$Q($E9QY~ � ��> x� 
 �?ǀ����JQE@@DQH$E�QQ~ � ��> x� 
 �?ǀ����JQE@@DQH$E�QQ             �                                            �          �JQE@@DQH$E�QQ| ���> ��  � �ǁ�� �JQE@@�Q|$EQQ| ���> �� � �ǁ�� �JQE@@�Q|$EQQ                                                          �          �JQE@@�Q|$EQQ� ���| ��    ������ (�2QEBAQEESQ� ���| ��    ������ (�2QEBAQEESQ                                                                       (�2QEBAQEESQx ���|��    ����� > �<"OD�<A�9�8��Qx ���|��    ����� > �<"OD�<A�9�8��Q                                                                       �<"OD�<A�9�8��Q  � �� �    ��� >       @         @   � �� �    ��� >       @         @                                                                              @         @    �   �      ?���  <    �  �    `    �    �   �      ?���  <    �  �    `    �                                                                           �  �    `    �     �    `       ~   |                          �    `       ~   |                                                                                                                                        x                                            x                                                                                                                                   >     �                                       >     �                                                                                                                                   <     �                                       <     �                                                                                                                                  |    �                                      |    �                                                                                                                                  x     �                                      x     �                                                                                                                                  �                                            �                                                                                                                                        �                                            �                                                                                                                                       �                                           �                                                                                                                                       �                                           �                                                                                                                                       �                                           �                                                                                                                                       ��                                           ��                                                                                                                                       ��                                           ��                                                                                                                                       �                                            �                                                                                                                                        �                                            �                                                                                                                                         �                                             �                                                                                                                         