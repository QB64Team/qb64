��h   2o o                                                                                                                                                                                                                                                                                                             �                          �                       ���          ��             �                       ���          ?���          @             ��         � ��        ����          �� �         > �@        ����        �����        > �         �          �����        ?�����        ��            �       �����~       ������          �        0 �� a       �������      ������       0    `�      ����       ?������      �������       �    `       ����       �������      �������                 �����      ������x      �������           �      � ��D      ���?���      �� ���        �8  @      �  ?�       ��  ���      ��  ?��        0  �        �   �      ��  ��      �   ��      �          p   �       �   ���      p   ���      �                 �            ��           ��                        �            ��           ��                        ��           �p           ��            �           �@           ��           ��             @            �$            ��            ��                          ~            �            �                         ?	            ?�            ?�                         ��           ��           ��                        �            ��           ��                        �            ��           ��                        �            ��           ��                        ��           �`           ��             �            ��            �p            ��             �            �@            ��            ��             @            |@            �            �             @            <             ?�            ?�                          >             ?�            ?�             $                        �            �                                     �            �                                     �            �                        �            �            �                         �            �            �                        �            �            �                         �            �            �                        Ā           ��           ��                       �            ��           ��                        �            ��           ��                       �            ��           ��           @           �            ��           ��            @           �@           ��           ��                        �            ��           ��                         �            ��            ��                        �            ��            ��                        �            ��            ��                        �             ��            ��                         �             ��            ��                         �             ��            ��                         �             ��            ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         o o ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  �����������  �����������  �����������  �����������  �����������  �����������  �����������  ����������    ���������    ���������    ���������    ���������    ���������    ���������    ���������    ��������     ��������     ��������     ��������     ��������     ��������     ��������     ��������     ��������      �������      �������      �������      �������      �������      �������      �������      �������      �������      �������      �������      �������      �������      �������      �������      �������  �  �������  �  �������  �  �������  �  ������� ��  ������� ��  ������� ��  ������� ��  ������� ���  ������� ���  ������� ���  ������� ���  �����������  ����������  ����������  ����������  ������������ ?������������ ?������������ ?������������ ?������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ����������������������������������������������������������������� ������������� ������������� ������������� ������������� ������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ?������������ ?������������ ?������������ ?������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ������������� ������������� ������������� ������������� ������������� ������������� ������������� ������������� ������������� ������������� ������������� ������������� ~������������ ~������������ ~������������ ~������������ ~������������ ~������������ ~������������ ~������������ ~������������ ~������������ ~������������ ~������������ >������������ >������������ >������������ >������������ >������������ >������������ >������������ >������������ >������������ >������������ >������������ >������������ >������������ >������������ >������������ >������������ >������������ >������������ >������������ >������������ >������������ >������������ >������������ >������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ������������ ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                    