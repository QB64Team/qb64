��`  �Lgm                �0                                          �0                                          �0                                          �0                                          �0      `                                 �0      `                                 �0      `                                 �0      `                                  0      `                                  0      `                                  0      `                                  0      `                                 3ǜ��pso�                               3ǜ��pso�                               3ǜ��pso�                               3ǜ��pso�                               ��l��m�3`clـ                              ��l��m�3`clـ                              ��l��m�3`clـ                              ��l��m�3`clـ                               ߷��m�3`cl߀                               ߷��m�3`cl߀                               ߷��m�3`cl߀                               ߷��m�3`cl߀                                                                                                                         �6�m�3`cl�                                                                                                                                                                      ٶl��m�3`a�ـ                                                                                                                                                                     �3ǌ�l�`1��6�                                                                                                                                                                               �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         �                                          �               >                                                                                                                     �               >                           �               >                            �                                           �                                          �               ��                          �               ��                          �               ݀                          	�               ��                          �               ��                          �               ��                          �              @                           �                                          �              @                          �              ��                                                                                                                 � �                                       p0              `                         �@�                                      p                                          �@�            4                          �`
�            6 6                        ܀ ��                                      �  �                      @ @              � �`            � �      p p              w��@            � �                       �  �            � �                         @            � �      � �              �� ��           �  �      � �              �� ��           �  �                       '  r`           � �                       "              �  �                     >  $>           � �     ��              >b  #>           � �                       ?�� ��           � �                       >   >           �  �      p p              Ŧ@Rр          3� �     ��              ��@R߀          3� �                       �߀ ��          ?� �                       ��  P��          3�  �                      �}  O.�          Æ 0�    ���             �}  O?�          Æ 0�                     9����@          �� ��                     8}  O@          À  �                     �D<��o�        Æ 0��     ���             s�<��1�         Æ 0��                     �}����/�        ?� �`                     rD<� �'         �  �`                    ��8� ���        Ç p��     ��             ��8� �@��        Ç p��                    ��������        ?� �                     ��8� � ��        �  �    ���            �8` �@        ?Ç p��    ��� �         w�8`@�@        ?Ç p��      �           ��������        0?� �                  �8@ �@        0�  �     �  �         ��8@A��        �Ä ���    ��� �         ��8  @��        �Ä ���     p             $������@        �?� ��                   $�8   �@        ��  ��   ����            @9  Np        À  ��`   �w��            w�8  !�        À  ��`    ���         �}�  ��       �?� � �      �            @8           �  � `    �  �         /�=@^ �@       Ô ��    ��� �          /�9@N1�        Ô ��      �         �9�� ���       �?� 	� �     p  �           8            �  �    �����          ��4� ���       8�H 	a�   �����          _�$� ��        8�H 	a�   ��          ��  g��       �?0 ~ �    p ��          \                 `     �  ��         ��R���@       x�* *A�    ��� ��          �����        x�: .A�      G�         ��@��       ?�<� � �     p  G�          �              8          ����8           ���@=��        8Ĥ ��   ��w�8          ��V@5_�        8�� ��   � ����         ��� Π�       ?�3 f �   �   8           �            8           �  ��         ��P\�        8ҕ T��    ��� �         ����_�        8ӝ \��     p  �         �� /��       ?�b # �                   �            8           ��x w�         ��� z���       JR %)    ��W�         ��� k���       Nr '9   �� xx�          ���h�       �1� � �        @           �     �                 �� �w�          ����
���       }�J��K�    ��^          �ߊ����       }�΀���   �� ���          �,}_�       ��1 F1��        @           �  �        �   �   ����w�          �N��.�       u�) JR�   �� y^          �.k��:q�       u�9 Ns�   �����          x�`Ǐ        �� 1�`�        @           `                @   �� �w�          g�GXq~�        Z���җ�    ��^          e��xQ��        [����   �� ���          z�>� �7�        �c c�        @           `�  2�        `      ����w�          �'@r\�         zҔ ��    �� y^          w�5�	�u�         ~󜀜�    �����          +8�09�j        1�c c�p        @           #  b         0�    �    �� �w�          
ϧ r��         �zR %/Z�    ��^          +��0S��         ��s g?ހ   �� ���          }��_        F1� �1        @            I  I          0       �� p           Γ� ��         =iH 	K^    �� yP          �����         ?y� 9�~    ����          �g  s�         �0 1�         @           �   �         @       �� �p           g����P         V�% R^�     ��P          ������         ^�= ^�    �� ���          >� x�          #� !�b         @            $�   �                  ��� �          �ˠ���         �� $��    �p x�          �ʠ���         �� '��    ����           �7@vq�         c c                      �   !�                  0 p ��          �����         +^J��=j     �� ��          ��h_��         /΀��z     0 p            C��|@         �1 F�                      A  A$             @    ��� �           ����׀         Y) JMx     p  �           �qPG_�         �9 N}�    ���             c����          0� 1�0                      a  @C             0     0 `             Z��ϭ@         ��AR��     ��             z�t^�@         ��As��     0 ` �           �ӈ�؀         ���a�                      �  D�           �   `�    ���              x����          ������     0               ~��
��          ������    ��� �           1����          c c`                      0�� ��             `     0 `              '|�+�r          {Ң��      ��              ^�.�          �����     0 `              ����           1�A�                       H� �`           1�  �      0 `              
����           �JA)Z�     ��              ����           ��A9ހ     0 `              s��           F1��1                         � �                     0 `              �u>�           =�QK�      ��              �]z�           ?����      0 `              ��#��           �"1�                       �@�           � �         ��          ^r'=P           V�"R�      �� ��          �R'5�           ^�"s�         �          9��            #��b         �           @                       ���          ����           􀗼      ��?����         ����           ����        ?��           ��݀           c c        ?��           ����           `       �����         ���           +R>%j      �������         ���           /s��z       ���          ���@           �>�       ���           ��             > @       ?�����          �h?�           x��x      ������          �h?�           ����       �����          o���            0��0       ��?���          l ;            0��0      ����o�p         \J=@           �b�      ����o�p         |9�?@           �~�      ��￟��          ��7Ȁ           ���      ��ϟ�`                        � `�      �������          ~�            ��      }�������          ~9�            ��      ���xp          7ƿ�            ��`      ���H0          6 �            `      ������          �r�           
06(      v������          ��~�           �>�      ������          G��            ?��      �����                        0        +�������          ��             �y��      k�������          ��            �y��      7������          ��(             ����      #�?�����          �(             �y��      ^��ۿ�,          �             ��@      ��ϛ��.          �             ��@      g�߿����          ��,            ����      F�����          $             ��@      ���ϝ��          ��              <      ������          ��              <       ��ߟ����          ��\            ����      ��Ϗ���          �@              0      ��w���          ��            �       ��w�7��          ��            �        ������l          ���            ����      ��g��$          ��            �       ����;���          #� 0            8       ����{���          #� 0            8       ��ϗ��v          ?���            ����     �����6          #�              8        ����~���          C�            0      ��������          C            0A      ���7���          }���            ߾��      ���6���          A                       ��������          ~8            ��      ��������          �             �"0     ���v���          C���            ?���     ���v���          B                        ��������         �
            ?� @�     ��������         �  
�           ?�  �     �������          ����            ��p     �������          �              @        ��އ'��d         T!�            uB!P     ��������         �             {@"p     ���"��&         _���           5����     �ڇ"��$                        1@        ����P         O�             ����       r�|`����         @           က�t     ��� �P         �����           ^�          �                           @         ݨh`Ĉ��         �9�            ���P      3_��?���          ���@           �t     ܠh`��         �~?x�           _����         �                           @         ������d          �	��           ���     �������         V5 �           �EcP         @          ����            �����           �                          �         �����D         ���            �	H`     ��������         X            �@Հp         @ (         ���            ��*�                                     �          �'�����         ���x            Ⱦ7�     ��������         �|�            �����                   ���             �>                        �               �        �g�����         ���            ��?�     �������         }_|            �w���          P         ����            �*                                                  <�O����         b#�            `�"?�     |�����X         �x            ��Aw�      �     �          ��             ��            �                                      ��� 0         _���            5�o       �����>�         ��G�            {��      N�\  �@          @�              �                                                    _�?��� `         ��            ;��       ��]����p         ���            ?���        �   �           �                                                                  = ��� �          ��             ?��       n�������         ���            =��                       #�              >          >                                          �����           ���             ��       &�������          ���             >��       ��                              @        ��                                           O               ��             ��       ���  �          ���             |        q���                           ��                                                    �&���            |�              ��       ������            ��             ��         :                 �                                                                                       ?�              ��                         �              ��                                                                                                                    �               ��                          �              ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ���  |x�     3ǀ   ? 0     �   � a��                                                                                                                                        �0  3f�       �l�          ټ     a��                                                                                                                                         �0  0f�       6`�    0       ��     3 �                                                                                                                                         �0x�0f�6��    6`��0�0m��    ��3 � 3 ��|                                                                                                                                       1�0͘|x6۰    6c��0�0m�`    �� ݀3 ��v                                                                                                                                       00��f�?�0    6`��0���`    ��3 ـ8��f                                                                                                                                       `0��f?�0    6`��0���`    ��3 ـ ��f                                                                                                                                       a�0͘3f��0    6l��p� �36`    ٌ� ـ �3f                                                                                                                                       `��x�|x�0    3ǀ��� �36`    �`ٰ �3f                                             